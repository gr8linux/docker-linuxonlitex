`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
m3f89l1Do6paww+DRMEVhGKd+j4DDOR84bBB8nJhTscTJgl1uiCl9jgTPqgBuSm+nURfqXjJo4sr
F0SFABDzpJgmBhgqpb5xopVntC/15p0EFKECClJkjZMrofmALtn6ap+t6jK1VH4UocirNIizxajx
5nCj+XIPy9KWYRfedaxEInL5yRFoKmEOeHbqaFWpyh7BMgYaGOGO+TFLodymMLtp36XHxi/uXbV3
WnXHUCyo2Tl195tba1qnP25Y7ZWIX4TJDEbAo45vP4V4B/dmHB4+OVIjaHHSkyIdVbZ7NdZyGeNk
/WlQS4KnkDTFagnPISFxmWlC3PLWs0H8uSjI+Q==

`protect encoding=(enctype="base64", line_length=76, bytes=314784)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
93FcZ/HK/CTqDgFLsZphTIWe0K2IgWtchd6KSgFiUGwcxJX+9/UKb/eTZ2qcUeMlcB5WSt1QuD2p
gjUthJedMOm5N8fT4Azoh2Zc1hpSJu18jR6wH5ILsnG0ktrk+47p+5WhxqPAXaWZ6ExD+yYdoo3O
W1Wn7PzDW+Yg1IHSD/+ZY3T6V8MKWKEfpKloe02A0Rpxf238e5BZyZb8GF3m4jx9KUlVmDRoLy43
X3mGFuWXn36AEm7K65l9+yOIpV4eCUoI+LiWWNmEf9HdWRBExnJXQE7TatGs4WrzFY4fOCe6nXR2
mVm/HfWyqkpZAHSdL6IuABhVafpynkslR9Xkj7vLCkzEOtxe5TqqhACfCLcXjvyz0zszo1SNOqOd
eoKoQ7nxuKHtT0RqjZTpnIdfCmceBaRDyFYKMHv3o2AMDgmFEojcnqeLOHibUoEdEdzG9d7L3c+I
drTQgtuaPCDQ3USMGMpUfG9VSrRSBjM+d/KwDejEYpDWI6rgsujMB4IeWCGB2t2bgR+EX3YaEKTn
WxtjpE2sqa+odR+Wk0rhLT6P/fCgKf6OQNXToVpM5GmOp6EarIpLuxC32FQ9At8DrF/H0sXke4o+
F0ZCF2wyaNKvvTaTG1X5sIDtWnYKiSNl/Ev1BGoFr8JH2K3JPHlF+1HIBO+jU0MZKY69aRmG5EQv
nO9+dgRacUlBJLhNVpMz+DPy0SnNIKRxNJofXF33TUSMV0lzkPI1HlKSSbwagbQRg8WPoWfHhAiS
Rz7A6hfKf32YkLRN/MWbw70vZL6PzOx9zHwLdB6hPtMTgKVPJd+861fvUzbiXHAYXBWRX6SNoVt2
0GBuH4iuE0Fq0pRpLfphETNQWLlNc+W4j/Vba1kmfp6Vv+Z3ik4uJwJ4WglD/95EhvqiA/CvkPOU
GH+m0oeWvpKVio7RyhQStOzkNSTTVPyKxj9vN12txFS18O/Sv7/FXTaCqmsvd+mPUkwA+OsyO+s+
DLYJnpZNdfZynWhuB0zHjnIM+wCWRBlnEpkQJBo7wbI70X0Dfoi2R1QFX4I4ldykhm56UEXIQcmW
doRlsVCwy0I2LBu+vIMrFH1Qc82h6BmmIEj5RQySTvuAx7KbNouRDAGhSU0Z3ZdNDCs/FqbXv0eS
fdJu06omXt3+wa6l+Ej8eS6b9iHdLheqyzlOERS+wpQlbWZoHWtd6Dor57GvlSCNqrYURAXm9SiY
ybgD/pleo75piGe0KU/9bKnf0RO7qBv1OQXQs7/3I1q4F4mi4RCqDkn/1011s/xoh7NIDVFsdJkY
br9zXW+di/XBCuPXzPWQibGN5kL9Tvm9iQbXt6wV6iRv4zKmEML69G6HVVJE6xmjjhrIuIsQmYDR
YxGKevipJJ/IPqgRMDbY+P3d2xu4HbfTPjhWeXfaUuFMlQYukhFv1+P1sjSBl2s97qf/6Qp+1P1p
Lpj0UCUwJm7Gs+XX7N4guQxRz9ULRmV7BGsp9k/2HvSY9/SOLzjpLvsstSH82Yl0IDL9vrA/HYOP
r8r3fYJqFoZz5QenIxO9WHpr4mc9sk2NJXzn1Z4vjzgOQ+GIuQ7wsABqI5/pDTk4cFEOeP8COWoP
hWFuvm1/FCpsHQXKHVDLm6H8kZvm8SN1+zatVJkXxxfgju0EmoIVFeLHPz6v5H8xmaC8favJrqTT
c54yFKsYXIrPgumLl61iBjKxQ+U3AJRxTHM+iWxNW1FXc0yVk7tXzdHq16qOmmC6eXPfVfKtEZk3
sDAGxahP9t0rdwrSlWNMtShGW2mqoKjB4Vd+oWLe8/qwH8yl0AGiHuoaMmsXdFRolu700zxoeS6v
Z+x7SxpZZeFILlX1wfM3aoqRx9zU84FxMdFabaQHCfxazJGliMRsEOaG5KcSccTlcXmKhyaabs/q
+Z4QTSvsDV6dP5vim0AcgVjYPKdGpH/x2CNvDaOOGeK9s7CwzimzEiRELZL2ayhSuP2djSpYqIO3
dtetREeYARTn7dY3LnNfXdiw+eRRPLfGoFcVDWM4+mSWbE7JgnVPcd/aFxeQKOK2BwjgxljnDVwU
KOKTaMQtBm6kJBMLbppxUH9LMj9NVD5wGzrCZ1NzT+0kE0v42pAPXrnzpcAk5Xa0OSXax0R/tkc+
lS0cvQ+zPj2ZjzuegjO8NoiQ/h/boGrxO8x9cJKXEAux+Yk0siKnzz5talTatnwHYVYoMwZaWH4k
O5NraTKCb9te5wZTVvusKiPimlvqHMY9lqHrsqer05F9NEvztLhF3qAhLmyQDT24DQcNgDlskzcc
o+JtnEQwgScTVJ8eHQA0JbiUlm9lTxhUa28UoqCmf00Cke+4NFEB7pkRm5lLPlHoC2shCzIdgQHi
qLaz0uRMrpbUBNhWMc9TAkYfQMgqHqIxwzvwem3BzcRhzBOooW3/v0ZrbzY4zwhOgjGVjDKF0zA2
sRDN45A6N8NcrP/e1B6TvAIwlSxggfGMamrJWT4m6trKariVys63ozteeR60S/bkSZ+HkIY3nZzl
e1geQk6HdsheaF1UQIpgA8XMpqOk/Sw8r4whFNk0z+kg4zXruIycKnlV41X2+6QsizYFZBQgHQ0z
+vDznIGel65PNCdGLNYXEn6VLowYfUPkh0NrJPBIbufIEbWl1q3I7haNV1QhG3WIzn6Fo1vANh1o
d1rJ2DeRSQyb2SQDbwKAsqUBf6K1TZupnNpaAdz8vXC9qw8dVfZsivlfeO4ymWZoapr1QeX+QTHP
YAYlljH1tpCz3Gzu0MsxEzKzck9nwQAarbgDj11ucEQOciwD09XmR7C0G4+q2c4Scpy+Uhux/P0n
bz3pMLYjraLzg75TbUD0DDo8wW4Nvqdm6fPWjq+4WyjiyhfO2l8rRYqI2wF0Gx2mW7OWNGqRPVfN
gjAO/2HHxAQQS1aZDaO8P54JnKzl1gPHkZLNjzgse7pVOp9OklSBUYAetIXzMHtTMZvOkmgEbpvv
9nPXXoSz+p+/7Fgiz8zh3AueeIkh5ha9Iy+IrUdWyL/eNCmyDZG8+6GAPVah6o4jRaKcZSNt0kTH
ecjzsdt+PTW4OqXiRK5x2+Q/Syg6XqKdbXRhmkkJEIV6eV0o3Z8+u8a4RwQA5DKgC/ZHlphCfHI5
oorltqCrbhF6/cN5sRFgput7rH0xXGYAUvaYKsFyKxJYaoEeyxc3geTr7XfGSCc1ynI8pPzjUNdX
Y6px6QSGbhMsQJJqIAG7g5SFVXFNSQ23I2i521SyJgbHNl3HOpFPNHDKgPjK3NP6lJcT6LpNpWMv
slIRtjiUZu0Zrs5NvLL4uTzHjdAjj7Vf9KnwZnBQh+BKjbHeLJqL3EUTTYZwCvCV9pZjVqwY1I1E
F8Bohffg8zJz1iVhNdphLIXFFx8wlQ4hdOTjzxqAkjgeCIrEni0yvhM9ZvTLa1xr9Wb4C1AuYe7F
NHIVSXaAXiqO9K/gMYAXJcAslguNUAhClLoQe8x4lpCG0/AjLglFawNGziN++UBMVJ6IRzcuIzV/
lvz9FkpY2eyQbVnMI6DB2mNBEBJloBzXkx/f8EC79tE4frOiXaVSZvdY7nTPM5MSxXy0o83pvPgQ
kkQZaO6pO9FcN31RIeaoLMQ38XXxPyY08jqUKlL+YGIdRnpFJcsJ8qKJSHclsw504UC+HC4hIlb+
Sovc5ivZJ9YsfTid3qUFngFzcjavhU7OvbQTrLwV7K2Ywbz/E6q+W5EBR2N+cHR2W1MmDJL/2ZNu
PIj2xUpua/6gwKraEli+57+jhkLYgdPpFhXWpNxZU6DkD4XOOvAa6/N/2bmLETYMmRNSUwA4jUxB
kMWMlKgXZojawJH/Z3HSwPUlH2Ntvs8wIN1+PNNc51i7vv/sPC1ZC7V/mNGakmx4pwla5vUIfnGH
4Mos7FH3yV4aRDZ8Fse9dtMibo+GRk2PRTtMa1jLv2QPooUff2cX3dp8IUgsqumDkR9uINQDtXkQ
AUZgGRmQM0wQNXSe2378ztEDyj7fUSD6BP88ghNVHs0wNeSDLzg+/ja6iHwzAAMaTYyAeEXEdiP4
S6iLIX0pQUKxadEsCFd3p32cL5iDfKxMkLA7eBymsmRscasuhz0V9kkW9NsYcmjHeZG9YIIVQHFR
P8ItNew6HMi41aDc0NdiFr+jAKJzT0isRpwjsFB5MTEWSHV1gWUMU6GcFUeDjgRhSyNyaSo+ipHJ
LllftrXUk0W8FsmTeTU/YUjAK2p+hy5GQ0ZHXJDfSntrZpko8TXXErO7t73VcRpUwaPfMtFBkn6n
Xei+1+R63dm9LsT0QBMQ/Y//vQf2M7hcVGa/V0l7aok3VWTLeSqN0/FbRwuGjId8i9MDlT8qLWNP
KkDNQU0MlkkggSUjUu6Jw65jSfD6YBPmIvxtsD/ZO5aUrgyGPjuMjaPgpC0FfChVsvFNg0vMulcu
PTkb5Q03u8KQDwunMYRnn9dOJ9ERAuEGyW2fbthx+PddXWS5shRBDjIPBvmI5JzMubKA8EpJCFUx
JdmuDJbweAN35Miv5mZK8wJxi/EBNrWY3Em7NT+3usplSCN6cdWAoZ288625hzMMuiiSW4qqcRiT
F0S4N64aYOoa6Oo9nRGPzajRuD7iFFkTkqv8TAY6Sy9VYA+fJhrPLCphg8r4iTnezGLqFeSVexVa
6UDKM+Ls4UeNh57nqJ8iNZnRLdKRGPCPa3ef+o2JbTo4h+3knzCtkwPqJ6FucPCZqSxEzh7AMw8z
r4zjnjQNg9MoLSPvP8CkknrHc4Pb4y66P9wpPavHFLkS7M6AeJ5RpAkv6DSvU47i0UW0DtZYCx52
7m9Y4l+OouRQ4cXaHtSgjnqIxRvTeSTrbQIjUkxL8LR1fxJsCpQbj6IyW8N6KQOfkVKsoosp2Vfc
ZC8eFWAetvKCdAXPsO274cvm0CiJ+L7ZAmhWCVGqtKr7KooRd4zFqTzXFN9QPTTp6ryvgCFmsahM
XHcEl1j5qDTe4BKBPWP3cjh1fp4RB9F4pmRU/jW212GTswTaiibnoaRVycbZ69hlJ0s8DHfAqFGm
HI49PiaNFCDM3pKiitmwv1+F13TD/x7Un1VzM3F/WerrkzIOz0Hh8pJTQKtqyfKdPNHgg5s9g2bI
EdMhChw8EGekxLJZ7NVqc2eLgyj4Ko5NufDSqVBg/PbIol/3VwEa/cyD18kxnzRWa0XWGmmkkmgy
F5rvquibYNOqfep+jXQlGjYpMi0Yem5JxH0nwmfyfD6vMelfIPLYSb5y2mZVpPjzLY7c+aKLVPTc
C6Qp1WnS6aGLpKdwyVhYHkZE2KTaLO6lfuU5DTC2EaVQcqxkO/XyAraN3/2Fa6MZeohgACP+kuw/
E0wUXs+5eF5VPwjBPQy5qGUrdgHfPD9xpt62N4zGKKcJa9hij561Q8AwCNLsGSJT0xZJ3HissaV8
gDcGbG62AlVnsGlTJMO1mVjSW9Z3RHrWJ5cMuLLAxB6wAJWe5uw/NxWpqHUFgpF5ZTjWYJrAk6sa
T4n/zwqWA2VkKMBdHfEhvWRJaIAo3h03BErA/bcK/ptoQNhq6WgzHC3vrDDBUrVOeIdPz4132g3x
H1EFGxCEFvo+0b8+3TFTo3C5rZlxxqYRjiX3zflheXnFaFxypSUzpUAcTCkTz1MLcwAc/dyDOi6x
SWNfOppQg6K1xsxoGrYFJucljxOH8KHEUKR+Wz9sEBn2euZn4xHdWeWq50MSnGIElwErFEAIaK+V
rGSJ2JlDSZUQ9rvzoUEKoN+MfwLYkOZ7ZTrof2UQr1zY4c6g4E2zq/y8/uJOTX2EcS+fDLwZgu0d
xfQcjQTJCav3BYWj3jXC4A+HkrrJFzfrtz/9Fd8n4ZWz8qGpxZHCMVELJZKMLNiE+Q0DTRXJRIwi
pqFLfKDijD6CXFOu533yBlHeLdiVn7/XtcPQVQr4DJOOneOpcSd4UVReaW7WLoNCnk1I1anKf6gu
ySVv8r2jNwkCAPDtRl0UW4HOzkrEu/k9kqV9conokTo/yS5Yxfd6SEEI91R2fqnnwkC8pIL/3Ldj
6gj4s4sM4bIOJRnBNYOfYjkyNw/c/ipAyPZ7MPwKJQ176qdWxNZVrqf2NT4z7wKw5qqBSdO82hPI
w1Zm8clW+ezeQwvIy8wzldYYr8nlYx7yqZ86UHSJ/fx6SAztgvV6UHRA7KWa1JJkDRUH4tC9zZff
DELR6RBXeUUvHvFvqpaBobjmMk4Eo8dT6mJ5PlJTOab0ccO4ALGNxzpVDY+2Z+vuxMd0og2/Q+gM
4VgHh8KySrTC53JZEvVP/cnA3F9ij7biZTSvd07FUhO2X5LJve12aTceo6SX7ltAXRTkFwMNEwI5
fT4eb4M+CS82gHw8fb/GYHyACGbm8SEeQLHWxfFJO/TFVIsEGTHLZAUkIse30s97qvL/VrpMatFi
wEe/IVgpCdmFb6YovQNUWL2J0bLmtU8ymUEmQmZbkiYUvZQU2ZssshpX5yv8lTfqnu3kbVSh52r6
VBOigNloZ9tUB1oOZrFF6MdRk4ay2tzDI/5Ax/HOJZTb3oLBJZTebI8ii8F/U42uRfBqyzJNWHz/
s1eR0w0fJa3A2Ch4ESWm48DA/z7+l4CxemP74VvZFIUVaNzcprkXmP1ziuYXTBENAxqgSCclJDU8
nhEpIBSUivIuDqqoyVxU6aL91Yc1MZ1K+4YdM/ahrvuZjhC+vkFo25a5nImasoQnXSd08RF/poTd
fUZFj/yDHpeuj8Kc4FNNcxmhLmUi1F6xrYuwQAjuM99UhaViPO9ToZc5spf5+0GP4mJIv8XVkmZO
PyaOtTQiht/Xjdwg0WOZHTpwI3kykX9c+5GR28dvhFzPEDE9qYGc4S9B131YuNJcHUiQ1dL6dHw8
1lvUddDp00ywlYdJCfWKwUPz+hStjGxwGcux4kwiumxr3vDm/iT0BTXE6q4bAiENP3MBgA5iHtk2
WftJT7XfJEP/TacwBUgx3bIOm1HCBIOlrcK8fk9Hl+PEwdl8XJoF/FLeDkxiLlFW1fhmVUa4nCSC
RLM5gibDCw/M2ah8FrDW6rC2pX7Oo/HRmfctOXmYHjK/Y4IwW5l6qGFjlGEkba0JKqt/TGBOgD6P
Gwg5Jqb8Lzei2BBM/BSaBAOjyVF5CpIZHpdIToMhGdzVQUXwdoy8d2oN+kb4rq5bkPjHMg+ko32d
Cby8NiHDcVGjVSnpwNcGHK7f/8+hRbM/s63lNlWBfp+y9w9HzNsBzj4JsRcmJKLiWAtDN+QUjVE9
kgGMJLDIMY7xkLj1iOao5RqluWK3h4D+/dUL8pOlpJBG0lEKUfFIFvUYrlvW8qPcdgnRmHSgv+2K
ZIGr/CyiXi7hpE7pDbfIG/ChNdZStApfTgGw6Ij4bYNv/kUPveRzjef9HkdZTbciJVW7Ie4uWdZk
5l7G3qIMJSswlX38PhLV6S7XnMgDPDfQT+d+ZPsm5+vcQAzxL7MZZWTkA+g/nf7Z9+tpVrC+AmRb
rV29CLaIKRm0cFa4oIdctyl9hCQ78Kcd4yFT+rUhzoaYcOTXa5fp1LH8cDCmDYVj9r96hbcGjWj2
tdZgQtUn6RH/dnsO4waF4R9FQS/RDiYk+9Xo0dV3t+bll1azUrc8/PTWBNYi4HBYhicAvsJT1KlH
EdB3HK4au2e7bxiwwyVssNv3uyb9qR3NxGCGZ5Jg6+s+uiR3iAPxj+Uml64wXQrrcc+aAyh81+Tu
UQe1Bngow9lOlrbKZ5zJfyNM28za1F8LgdCEsYdrZvSm/IHTFLP8ropnABYCUcCCsBkQIPKFt/vv
p5wgkw6bUfzG0gqn6kNXx6pxpLmuJGS0giFB85ujTgserd7WWw0MYd2N47/u/i9AVTUhbxvm2p6H
TGvl0dLToIx2ICMaVoenYeJ2McFcQMlCITi1F4Duw058rDGDod44E5dbZslAxhjpxDQicfrB57dH
AxN++fyJuVvYfnupBg79UuomR6csEYqt6MCfbsux8W7u/lcXGoqS99jKBZXiGkjSH876imD7xvU9
Vb8OQyHDASISHyqMWkNcXkeeXWQhaEs8G/EQ4KjwX3ucYuTgGhEu1sgHTV6bXCiSRpMM4VgfHgx5
mwawKQ5ElmN91JqZQfqBdNQkRyXH5J05T+g4rtjv5J8jpWGaG9gf3JYulaIJ3jdwDPAYDXmVJeEh
Wt7XfmKYF/8fUKyNXOJBSewiwdjMfkdSPyldw7HsdWcGxfmMwsZGP+rsJZ8lTIMna1KJv/mI2dou
IcjzyyxDxVZV3OdNxq1NEOKeUt66VD35XhWYxDi866mOZUKkhFcXuazH2hR2mLJ4LAAfrPtYEmfw
7eaozQiGa8qT0yZveI+ahYL/vmOmnbz7TsG+pdIbe3/acg4F9zMjcNh1t8Ro9zBIdoz1usxTJ6L6
ECtNEPMQAL37zRyn4Py2f61AE+NJ2oo9ARxqCXU32XMvr6FTiuBGpUH0llBysflFbLnDhrTGeCXE
9FGq9FYrN2U6HElsHTCO0x+5OQISHJVl6ErZDDWTm0rkOV2BxevtFEFX8HyEkqz0SmCIyZkg50m/
pz8SD3DnNdmsa8Tkq2jGBT54ic5F3RWHXvq5WO17hfrsalPxPdu+kM5Tjs9UowQX6+anfDZeCzfw
Gvn6gBy4zy0IP3IUWOP35eGGgDlZHf81UWKASa0Fv8auRh8GBZxftfVp5KSokGxbxvJ5Jp71xTSS
u4/U7yMklhp+rfa6mt3B/WUdfQfl1wBjUkM005kCRFUwnaj8tIDQTvWCB2W3LKvB3THtB65cUr8m
1h6szhZfise+tFRsXL4rHCogkuIU9CkMkveNoXu+3dhYYKX+9YOIfzkoLCyThgeFZkgPfL1rzzxo
AhYBIzG9z2LntdWEmrdH5wlCAUfMUduWoWin4KN+7MUeA7hWE5xy4ryzIDxlZZ5TUcnYbIqXTs9j
L+hFNOAwq7ifyxeBdlrlLRwCYELTLZt9y5ROdUTaixMM4AColWmn9+ywGCSVkiwCmOIUWiQsDwJ7
IpLx2NCPv/kZEgFI46XYG7xICCC0nalarOE52UKdMFCP0fNO6HB+z8pVVCJeBL9xUtl+QgxSEcMM
K7f42mS3ys05iM8fJumIpst8Lz3/5BvJWOs6Qgo+DTveSLN/pKNdVcPlzPQMZDouPBLaPsiAsAF0
e4R0qXrL1KAYDyeBz8K26DR96V/DBl5ZRJ9xvNugwsyvd1d34NPwoZZ70RIEliQfCyWtioQK2uA/
NqaX8iKwBif5QpBgrD+8ukb2b4ZNhkQPL6jO7p0arAWrAUz0qgfRXY8T9NVzFtORMm4o1/dtKjjo
hoONpI0MQ3S7ZsMPAwtszgQTAJpHeAE+b0I7avWTeF5UT8p4bcUPRsGVKYQDB30WZnV1AOwT5zWu
Wg3iTs5B9bzbLhvCJj16wHmZO3SPuh4lwZxivzE8oTrqdbRVfJlTFUL+YHRroKCZKhSoihtXSw7C
OC8yc01iqGuAAwkU8WThPqzVmUyvtmpdjk4IjRYAjDYHptSNcFHm7jPjpH6viKt25OTXxSvve4NW
rGF+bxYUa9rRFagykGcUa+/cg76yc7SfVrBplQQgV7z+Be9woavVjJ+vv6QzNAjxoXX9cbwJ1sIs
Ox4mZ8Avcsyq3ElyDRm6QuHO4D8Vqtz0p5YKKAkHDyfm52U6PJNvU/xBhbMab7pi+6k/0O7/y5fl
IPTKB245viOL8D95KV8V4ks46Gnhv423M+preekuD7hfMtfiWimliWAsVQ/M2gfJe1cWKpEkjMEG
KapfGt38VgusvjEXo27ukP+tzjdoaeR5GUlrHya3Sww7pyUcgXuQFwj4stvL8PktGPo9ksau8OGQ
zEPv6qr7c+xCSl9MzvLe+CyVj6ax5HFxqSMJ5DBX5i7l1vLLfHJRUng8HJkMk8Vg/U52rlFoQW0+
cqe4TEcHX2e9AEwpVKF9uNzZBSI1IqRJXB2qzGb/RNWv1HxAW3QlVCJaR4H9RbZTCojlzsjFTjQa
A4ipAxpEofBTkEX/QReqLvX4QLvDRox8HopjFSScFnyfaKureYthAFfVIRhUgNRXAITBXw32zYss
36Ackakfm2CqDSlgVBDYHXUYIrFaF8fsoSjuf+awaBV/PtaTVS/P0Ar6+DSQNi+eFgaTuYoohQBU
QOACAGEvOZJoxKC0i86fX3FCG6DorvDJTaaVlujLcXo0O797Ex0kMrKTEX5ra9fus8e6Jor+DQos
eyBSQVpplE2utIE7Nwv3DimhqjfUlCJI+nZw+hdEIgeByNDhwzG5wMd8+doeAfKdNKLL1+HyewL/
v9FPlN9XvEf8dCZ9cJPjXKRfbc8BIR3g1UhBdYHF+Vo52NmLOn8Ri7Mwrm6V0IlbsUMQqogwNYzQ
z40RtyaInT9zqmX5TvQhUIUYRUVpWZEM9+yWTh+6woESk1JboQbDFkkWRglme33bDniCdSyZi740
Mb1cNQo2Az5DnH1m5Xe43/41Ly5AZL+LHH93keMui2b89BfKmeQZxQEi64RRPJ5solPuqnejGNip
WTjgvyBgZBmRKe6f1P3f2n/zp9kFVnwXpflBHjCg1wWBHpqdjl2+DZyhW7B8gB3K69Umm1Bwmqm9
PrYxR5ozildJQfLEg/+7tte0GNxgfh5luixSjMvGQaoZxYIdUy2Y5h7EpCSeKojZx9wbVcVuK3i3
4+4T2cxwWhkzTZefby5cbNpL6YisDcMl9VxM/+I5Uw8neHwnbKgAAzc+Bt+v246Prk8goksyBagV
ReG0UypDQcxRofvwycEV3UA5Pot6yrIki1IJM+okt2lbmdw7vrXFWcFacyGmfJ3AJUd9i6iF7bV8
0haeYeWUIo6rosEXkplpafrtoan4mQRs12CYG1XajlEppKWyYPajMoee9Ou01Etw9t8aa88rHPvY
iJuCqbUlbl6WIk0HZLG19UYIERafIXKYcsBgirLlc+Gypul4OC4F/68uA0gMgbvMfEKQDVZEiaLr
efcOnCaN7F/nMH2lvORiJ3eswnUhfwUwR1Q/V+HiVV+PyJ6pe9v4opbxviVd5/hH00WGLBdoR1Un
n4/2dnTkAQXZKZk8WLNU1I5bo2YNXxzUy3LNvOD/mroCDH0unTxEpNgFg3jbUiNtPlrzW5VtA5YM
hSKR1u6nUAnLcYGC4GU5q0N0/k8sUzEmPEafl5ZeiRbAFE4YxT+fE5BbmVP20E0UZi9Y86qoiOIU
qpcAYZormQbv+wdZ7pnTn26717KHrPEi1YEwyYuHlEJWzcEdPeiSeHraF5th7zS9NlxCcOxg47+0
2/hJM4VIT9L/oKJmtI4Ds7ldsPyWB0MOJmngwDQG3hs+V0MloFYUQpmu8iBn61sAhNvG0ZX4daIl
czuCIX+WFK6hvDVuFbPQG/YCWguEjWwsljr+P+6d+bfWuagDqPo6B7bKjwf0N96r0gof2gOzncoq
xTY+x2HzfiODRYRs5rV0bP1h76tnfvDVlV1hm0grQUyWuDc/PzMEz/ks32qcjaZgLyf5rT1UNI4T
Akq2bcU8GsrbDKuYEsCNqwerBZ0EGWS9tgzpdUOognDUOVKmHEwMG3snfrseSuMD9GMUfMsmxqsz
yhRqeo5SxHEszTjLPEvrPlA9e+JNAxUv8hcrLPVlApTDiVj7gFTHnGRUIaakOPeCx+Aq8r4Tovbh
4ttoBQ7Qf65ju6PnNWoizBgM7XgaO4DuSbl8osVrkBGLOxPh6Otn+57GD/OzwrM6s0u9tGw/FgAg
PV5V6r3/XO3dyL+mMllRnY5kkJf24rjBArm3Z9Tr27pZT7LZEXBptQy6qmr38FoI2LpdwXmVEZj3
rvH4e38M4pGlNvv/MpQJFAKhDra7w+O9zs5DrKbMQ7pieU20CjH6SWlvFWSVBKapCdZqBPfuPww/
GNWurfxcUiXC93hsIoighqvMpw7zPypU8S6zFuolXEwJ9PGY2fXyNQ8miZE8ARfLboBLXyeiNmL5
gICOtosSSGcCaLhBJXv9LpyW22KHzxL+oxArmIwJSmf+KC/cs9t8F/ykweK38A3upUa0IodzMJss
3Vq10FAnMk7avAZSKtvLJmkVFV1AEkt2OSfYR2LEtKmlLx8jyJoDqcNaUeDpUtPAITc7j1kA8oJ4
pnuUW/SW2OO1erw6BeZbcvLFe0EEMYKFrxEDGX5OjL/FdFVxLsMXBuDLJtY18RsS1sMi5G0p6iUt
6W+eU6jCmL8K+pSE52HC3CiIB/GCk2IezIlEsvXTMGFCKsRZH285ttoCMdMBGGJCw2d5ZUPOzqbi
wNqnKaXIMudUY213U6Rj9OoH7PYfqlmBEYJXG8T25wYuREdsMLL4y0eQqN6esMDQUg6ms9NcuQJy
duUhASU/2XdEvvEkQSe/XA1xzkCxm6e1AR7BkXN6YlC4jWNEO0QQCV3nCPmZIdPXWiw0tPdM9AUA
p+7ZcRi75HSvmhctBrA+ucHCbC1g/pkErgUPhxTqegpk/qz5q8HsKUwC+cakEQy9t+FTkj9MlGBY
jvTMNDIMiB/boSa0GuAxDhrN18cyKoaaAXsQQzjCeU1RXOAI3Va+xtRJB+YaBsvc2hTwcNI9uPP1
2oKJsu+HwOkONrljhqi1fUBlcyF5XbRQu9dBKXJHrvhabBnq7iFrhgK6UReaoaygLkKHr0qBI5Hz
T1W6HOY373ZhFuy1Jv9dgOogpE8wvHrMHDc7ZMgUp0EI0fE5X5s+PDIpRmsokTHVixU5ERzUMplv
+2IEZF3HfhvHLdQ1dh6FVBlmFCoyqYHRTEDFPHDdn9tW6n9pVLs+vbIhzGv/pfvDfNA0wZNI3M90
J5tJOb8ySyKfpgDl8kpyeRcR2QpZm6C7Ju1tfAlNJ3yGeJQ4r0Bwfadx3TdD8ADoSnSpIrDNGFIe
KGpXtLo+Zd5MvdZ/MQHZ4Cbqun+6mp1cCYI3btpuh3XxBsBtQP833mnLoRO/FjNqbjjidWiykLFK
sNZfAVJ41GiCUTd4nbxEdLEK5YON0CLQxqN0tHqoS3M1bLb1At5T8hTxkAXmHCwj8rGagdOQliOa
pUEbHzo6kcSSdOjVF+2inSOsscbnOrLoHWe7AGtF+eMQ5iqo4K5JsWO45RzlxBdRQmQZAQFhAcG2
jYuU1MCth8tciihNFUiSWZi12rt2S+bWc+tR9dGmSiF4oyrWy9XnrHjI6CWnVuT/eZJsUWvVOCxF
+q/tD++3I8UIbaNvh4RQn8+ZamcWbujxm+wXbCPU//tqCO+BD+LnnDtLlaltTIMX0gWe8BahmxNf
E4biFQGAUFxagh4pOhlbfQsvIg9e3mJpE0xxjNOWGC6i48djvDmlRVcQ9GTcg/Uu3nRwQWwCc6wo
Mr88AK+GOTK1VkReDKc1lQHIt+CqFuFX0lP5HMMSFkTwgyyzI8AHKx/++QWcWw6zcRXAKEP/XsF2
zSTqe6iUTattTHSbbhPrN1ryaTtwl2raa8MfEqlSgThMBeo4Hplp9Ixb3LxBohmNsyDX26cYSt6R
+OYl3erLe6vAnqlbU1NQ+9J6NtTvWtsHk2Aq6qbgTupqw5NKF4hsXPefn2aCEsTyfXOHsjfM2P2m
aJXtbHa5Qn6HSUWMZFpXLumjbUCJA9pWcGxxqgZ7vh1LRJtnYHUP/QhPZPXrh3WBLkLFgYK3HwV5
y3HZjJ1AbiQKOEV6lh8RYww3Z4MSMdx0d/5xfD4e2uJfUSsGrn2EmB6e1sx+VXs4fMzpFb+SAdq+
Z74QXBGivg13MVbQB9Vjv5ccBhYVhVw6n2H+68uBMb0QLauUsk32MtLbwtfcBWPhphhkSnBLbtcI
LyuztGqMs3CqIjhNx2WBItBTgYyDr5+sBWNZVKPBPfx+gJ71jFakmndHyblOTJruePeA0tjg+9Oe
8Zdkl/43i9uzmf0134rg+F+6bQ0bMZg3oWAhvLe4e+1uAefoldcPTp2A2zGNFTtdOUGebmZsak62
jUY421yFeLiptam66vlVMmn+90miWf/QoUpafBcI6w6Lcs+sgFDXjy3YI2WJby62FwiU8iUBxGav
1kAVKoZSryzYm0s/nOYceG/E+CcFn3ojrbmllb6wg+EJXepEdbMcVi99w/OUju8S/pKPZ8UnJYaA
gWYkA5RbKItDh6Z0WdV0F/PBzYXJS7/TmvxQERS138mziSCgb0w0X8JrNgABOTspwuR3U6Y9NPOo
5Ys1pF+GyRJo3fcOq9lBkk9GjvUoErsW+6ay097uBFyZyunFdm8iAZpZ+86HmIeIpNVd1iTO3oTa
WNoneev4t8wLoD1UhEw1mQAIlrs9KiaslpK1xVuz9XdFVE43lNEygvLObUuDuD770ozKH5JbhejR
toX+WV8fIEw1+nUbZtqB1xCtpfuGv9RYcrG75Nr8Jl3FYLFkMdgMk/gXgHX0cLcfQbbixgBuwTTK
we4OBPdT3HL3Wpyt843yrj0c3u85yFEO3iqhzvFfrUuWC2wFH2QuCpEZvhzRQa82ws4AbLpk12Pk
1QJtX2vZbStecDk5cqpFaACdjUatWgN1JQF0z1PhTzyCk0UIMdpCGkbdj7TyjqIAO6gddxPzQLiX
vahqFxSdETYa20MMrHoyM5nmdrRxeMkRLYA0FXePFkWrlIVi0VrAO9JqbYJHwwlMZW1bgVbxJjUr
LZL69lZPsddY8//XKC8QbJrgBZvhtQbF/pAJjqFgORsVYnA1jGR7+VN6/ZDjbCvxtmbSX0bokGTp
6WtTDFRPLQh1QLp4dkdj38KcamJI4IFy0r9sW2Ww3imSrcfKj+c8QIBiZQ6kSrrHR7IUHmqorjef
kPLco1zKo4NEMfuNmZlH6mMSuQABeTgp1adYWZhhHtwwDahivGpQbsmVxNYB67A148ImjIFLRNit
Z6K4hqUsbX+uiyT6ub9QSZt7Kt0XLICV11PGMaCc91LufeBbad22X1Of6g2RlaxVwGqVsvbkDoEt
FIAjHfXa4YZelPmBA/rWX+oSa+luPHw9zk796QScyBhROh1tbMwFifNRU4AEUl5FT8uxupRede7M
pw7BYsrPjJx3tKSOs5OGdcbCpccUC3wfk3tdQcRFDwn9fXwQZo2wAeruonJyzAt0KswY219VLMMQ
wEQT6tfzk7JOZ14RCUdcouDNcgFg6CSmkwYIL0rJGveQcE9LgGYsvnqP1Tvv186nsnYS/Y6MeU8N
Mul4IdZszSH08Hn+qA1fjqtneds0NkEiDq/jACb0lfqEfD/skKimJVSO3YuPSbODnYW4kqFKJSnr
ScK/aKony2S9JfE1lZYdgZ+yotBh6LBpAMxZsKVeCx5PKb7M9XzG6gWQ8LxUJ7O/inktNV6HXzou
wDGLOMyQSoH/KWQShy4602kxJucfF+DhHv5KpAUgC7AC9xXvAfn1RBKRtLew31eSzPn9FSxriwrQ
fWMvU2iR+f11LqwULgaHwqnAvpHn8w56SBo1ThaisLz4TPm6lsY++YbkAq28dQJkIEU2NPg258Ic
phtJBKtWRZ41oYRP67/2IIyZkJ5g5XcJ4emFcYy2p66OxRCmVnMTYuZiKgpv4A98H1dVfUzJJvoo
31jEAAknMmTFVmETPWunrDIDeANj+QxfjWqCMm/mZg1wCkaGNXOa8mw4Qg1n5vH3jvF9577ssNrx
Ke1k7VZqyI7SJJD2UQzMZoQNAodjKZ6gYnTfKK5T1t96L/MNN8Vi/cK4OBSvfNBGwMSFUl/WIcZF
4ePnr00eGa401qgAfXd8vkNPmjycj6H8ZSl1k5NSnMcdVFUsN/nkzrL8RfkkP09k+OERzhHEGVi7
jSVTkVadAjf4UFrvuy7wIZJG2xqafzkmNBwOoR4b5vVXi6E+a35Mr1otMzSikgtDztZoXuwRQ54i
olRuUqotV+57QBdqqP1FXiDAne62At4oVm2CtcghtMHZm2s51MLqJ2BC4b3aP7T0jB7y6pphs9Q/
ZTrp8IvQ9Y+ZUXm+6Gf0v1cRdd62XiSmUFlPuJpikyvCkIXfeQwsysF+P2ZfauuRu8jHXOFLloGo
Shw1i+eipVBJzBI/XSrpavhCdKRpHrbyF8xxcLgymNzwxrL3/LdmIw7ohgEKf3KalKfhCrHK7M8P
55QK7d7adBfZ5IRDt4qjo7k8S4buD0C6YOAb18muPqiOsrqOhKDgnol8tBFOzKwa9EKY3aF0sRg2
o2Lq19yo9bKK4BBkhhlCLMS2X+jGff5mWoSEnYEobeFr7GJPebBDpKZe+8WDd7pC4ZAvk3wuyzg9
8WxUb6M64FkVTC9TTcOQrOUuAiIXrA8Ioc/NUF0lF24/VUOq4IheCA6qy8DLNFiNMtJCduOxko1V
Uyue5wmE9UQPwpC91S+xBXPF2Z7KLopJizzZ0DrqEAqmScBlywPGDVum6NyOH/QYvST3072Y2bv8
OH3BnnqsJ1/IHmUG7bxbOZ4W8Qygq6UOELO/YnnjWxEhjZkrNCuwjketjBFVneEZULooYo/7RwhP
HBGCc7LlotYhDyMkVVr9fvzOIFEHv3SYJDp/5QPgUr6Fxifs34cXsu3tO+UYTjl3oHIXwUijkzaV
OY5iHegdg8/SvPI1uiqKlkHqaZ1jHGnxgkUyYuQ1t5TQtlhEElUQ2CMVRm9xAH46VxIQPQ9il9Lb
6227X9YnedWQQTjA6zX82ONdlnZrCr+JJ53fDnGcTHDhg8WORdHq5YxRjQYTICP9Zik8DiHAa3Me
4o48eog0GQCiGxynxFSLc3DpUnRpIn/BUcKxo/8FTEVe4MNhCvXxerjYNapNFPa5CqI7GaYeqfJE
1Pr4dHIxtdN81sdQ76bkBDuiKs5xfUzRFbRV3Ellr8I67KZOAExFmAxPbXnipySxAOhNg6qJ760q
mQrUhfw3Je5ON4pxEb5812ubez8CeI/Qe5zjkdE3mwcE6AexJOCHCW1/kcnzHpJ2/VfiOJ6GLOD8
XC0IcIO/9jNucydu4mjiGDQICcYSPV8cjwZtb9S16zd9mhxfL8dFEp/PGInlt1XqS3PIzS58kMXR
fnytiV3dmOlhEnDqx01XxWNdZ7OeoCnvdUl/qC26g+gVC/dYLWtmBkY9iPK7GW1buCLjCAU5+KIb
wTfGEakNjeQVhqlzph1MQuCu2FlSOpX9Y5A7huQVVHwpusfpDmZ3esNekR4oxxPRnUNWvyAdeDkD
Ynk7m3LO2irHYMI+eucvTuVsoCpq4nv4yqBMSExewG6hpngKvik4zTinU2uIXkgKSX17/cgqKK0x
sUMIaqoiN5uhvYXwuWmAFpeOuwHakQ4CbqI1xKaIbrRVZABVKq9oeajj25e/5Xbmpy85uHGCNfL6
XryqZNuEhxqsry+vsWmkE8TL4Iskck1bgo+iAk1gTsnMVG4s3AneObi3G5M/ZKr0FJz0C/MlQWaA
d9djviZ4QsiWu/2VdNJhCGVesUPaVT1N8SV1w780yELdBNlTsOGSX/ADHyta15RO/okqXEZadequ
hVhAqPdZDMqMfAgczDxrASDCdOyoq24d2P+DGcTsN16tEeigR+fmPPR2WA+kt7twoZ39OBUGMVfy
+553iN6lRCfcOytNJE0Fg85rclBaNaF5mm8JMMO/ZPfn/cNCJ2kwu4ZQ8b3Z1lR0LMVrglKbHD5a
M7utmBBU8E7/d/8dBggVQfwFqlNIUBU7C51PWs489qADTGSG09NyiVkz1lyUQrQCC+e1UyQiSGB1
C9WDN3cGDQOL+pIdWS4va4b1db2VmGfVmF2x4wyII0zvfOaaRpNw5EzG4foT3l3qtw7RODlIXbK7
FlaDbnsA7ZkOqdP9CxC13oIghHDlm3RiIIZYXXwawQgLDbNMLaIQVszJCGSGaLsamUjdWDKqgKm8
ftL9oRDvbR/IZ+st1M3w3HY87UkhiL5mo7vULTDb4g5+x9FDdAYS6d1p5faqfAqK6EEJ1GVtXxyp
3HFM9QVo3XpDjYXJS0qQEAY6+qLV/LorePblObPfP/v2lI/7ca3Ml3BDyRvF4/Mf070tVyZuY4Iz
bbtBTJshtGzNK9oDc0H1WhrSQU/A6Jgh4eWyZfU2Q7IdWjcDSwUSYADQfmdxzK1jRwn2yAkQ0/sv
oH5a1sovpPTYTjvlJqzdqwgmVrFejgaE6wlZ3vCNmObWueTkMDaSck3Lb1SJ1zA8+pDH3vCPTNMK
QlwwLBKaDjPWvIAsNcfPhPx1aH9bTycOF5AHvL92HC/mkVyefI7AZfRHIK9HLykSmUnZmBdGFoAb
lOCpNMdlJaxlSriQ0GzwQrb8Z3mMonmYCh2tzO3lYdBCOLFSAlzcEKXWZcrbZiF9x3rWUlqlJjEA
U880LEpllF79CscRX0/o7xJbQ6e757EkvnykzphvOT85wFAzZDdx0crGK2PLLMm7c460dudieeT0
2uniaizwZ4/WnuETE+h6D9cf7rsWAR74ceMHuFVR9l2eH6G7TT1GErMwV/6XLBKDKVpNeGC8AwdL
CXUNwNUSJbPPzFTlIGH3piGQIorLC12iVkWFibAhQ5RUUtt4i3XmI+LoHoohg4qOQ9+zWK96pwKD
Z8jU5E/hoPTOJkqev/RsM/rD6sNP21zAuzMJBd9n9tXyuYrFyP22RofqYT9Kdit77XAIeOuzJozJ
N8aA3AzqVbpblDfnbkbo5EGNvWRb2CRIqqM6s+GLArUnWdK218UBqAbrbeXik4idxaASH+o2HQUj
GuT7xBQjWe+w3GwXQUbaQeQD10m3cyCLZyn67mMJyt99FUwWGYkiDK4uICA7DEnMAxydR4HSkhho
YdVTduFsTeclZtnHHBOdEgixUO6MZ7M+LCoFJ6Rjr9IZPz/k0zxe6LYPawVmepP2+47/09VvGc/6
q5yTyvF0TgRZQ1uPtOgm+ti9YyO7GuCMYWl95Fxg6QdbljAxJ9tKkiBndpPmCXEtkm3EYd4oI0aL
XplTyS32LP9ouxErr1uoE/q4EIIxjpKaf7eGLjZum3h/dwvO0vOzlc7v6G5bFuN6NDCsymtsWWOu
488pwpGHKCEIG5NomVB1XGaZLN8cDUrp0rtNU5opcY76QOYEZzOitzjhWJX2SBSZjePTes3QW3CP
7TEy9H8xCxLYZJ66204AeFJJLZlHNLLuOttmZWleh9giTpP2H7YqmbdpBy2k4ySEqZHldR1avT2u
DXE0929yFJ/nh6/IvAVRZDQ9ZSzBVl4K8ivuPVt0QKW+KlN0ULpZqMveo+XrVeQjexzYYjF/bTxf
I1C2phf3zCU6ILEudgVIgT3llCgSQraq8OVAfE490Ke21xhEd7hw+btGFR6qHu5+kp8ES+sFVZuI
uaH3corq5EC3buMx8ugYUdrNix/lTjHD16S7sVT+lCbFmgXO5ZB9/qzfQQGBzG0ygcM7MBZEU6pJ
iMCm6Prf/xcnLWv/m7aGSm1e54BUspVD0UB+n0rxdjMbCVro9hHTsXNGLfi0os5OnpI4kGoKty0Q
c8fETPHPRTsNlOnmBssWE20ubAEIy1rWvbcSntKw0J2H6Kk8rcKPqQjwvPH4UkgIiQ+wUvDNUnzU
pN+rSL7Nbp3KmK+RlsDweGSSe0kA2ylBl/Dp6mET0SEDqBo2u3ALFz3nTDh3ZPdwFfcyZhHlCXJa
LIWXt/59C6O77GibcQaP0l/YWpNEqdk0RiiZpUjglqzH00mtJG9Cf6eibDABnf13Q7qGCmx2MCWq
2mPC2d8mk65qYtigdUpOMRnAglB52rq0hOQlcyFNwmmKUbxSz+yZawJ1wv7S3qDKtpKz4TWUzhbc
N0obTnZoPQhUmoeGVw+Yaz9CGKSBrzvJ5meEPX4pw2fnG4xBhb8m43DWQFDJKvyAR6emMNSz9IeG
Bk40NjQ/3zw81GyNfKq3EXlKQqXh88VEEDoxLOdbhU46eEaXXd93BkGMDKZ0LRqRaPo9bYiIxCjj
GOP7LHDEipudD9f65jxLnkPSELScQE8t434V2k0Gqco4Cc4gIKMPzAJ03x5FFmCPUAQahn3td3yH
OcAz+GKX7Emb/MoGYhH2Sw/iFp7ryrXp2h2kA+BBjifTWUwJstp0vw6CnqaW41uq+R1EpWMAR5u/
ZwPN2htRncDXTzzhwzAEuf8yK7egxSlMkV2bHlZsLexclsgrMvHrcc8//g0fyR/xxBd3lS/WeNhO
Qcn0Ziy+cVgRRJjt9R5+7pHF393K7NfyHIeySv0TAe+MBLrAZVI17J4t5LxngKjiEzBgKPzFc1iB
b+mVt3Y6eTWS9+SfH7yZyIIpjSFU5+NuuRXXoDmqgswLh1ckskthZR28T2ANE/LvM9orvZ/7xmCY
TMSF60XFlIyizyHLbH+SkSPk26Oo6Eldva2ngc15QwGsUDDT4PsnFW3+wUDxxSM/fsamdzDdK2XP
u/M3k2m5qq6vVurr4Dv0syiah98xUe0RnRC/+fKkRx+s48zgb5OkgCxo6KD+qXD/m5G6QwCOC1Cs
dmC3nRLMoVNWobjs3omz0KGuxLVpYOEqt62vfwauWTDS2WVuvKJAVmeJFWWgpQ0YQ3H/YowiV2OJ
3PWJYEOUvs61PYMtG9rnMXwPc4ltqSdpbUj/azQG0KVqhMPDwNzdNlLLV31QKrofxUx1UavGNoub
/o5SgCA1POJLgDHfhMBfdyG38sdJskAUUvdQ7SJhaswFop2gNwLvbZD9QF4++1B3uHg2FDRcieUv
k4RIk9BTAWjH/tX/heCQ4CS8DqTJ+YCxgmnSJlcNROc6PmTCf0UfHHMD3KXh+G2DqJus323alR11
1hPu6pL5a7f64LKND9kLitR6Ee0aBjoDHhxTMhATqkGQU3gni5JDxeP2gKP4RA3AwbHxRtl/4SEP
HmcFZ12d0Q1qo2TFE74Nd3YrZmsSHqqGWTOs/ta+WSmaEZueVziPZUmnxxVcSAy2q5o9ejAsReHJ
3reHn8Tb/i8rfmMSYw0Tc5gIzzqg9JiqrJxH0epfYPUDt8t5xGDnKGNgXJFb9wRZuswgqije4d7d
8ObNyODCneEH/kVwZshJC275CFe03NjOem/MR0e8k8q8/x6TKhdcyB0CX122G53ZCaQRF+Ff2rpV
7l1iDZpCVjMadEydkEg08MKcPj86+T2XAaRM4QREamf2Vt57MqQN77WWjYxYxp9FT5K61cHGAD3N
YXEkvie7nC5CyKDCHBZa13u9DE6nrh9zBi4hLMmuT7RMfVc8GFWc8LaYT2aLNkA5Oj7EyvsudyZZ
bD2d1ByOWO4F/Ia/5IN+iHgFCiThLdjn8cTeedDfOGvnjhVJVWoJwR/1kS9I/1Rb4UlrZ8r5JaZI
77LWnTqN4Ge7RlERKcbSB0660cZRnDCNHvzDguFEQ5lePr+WdsDKroDsLLcvJ9npu/lklP3x8vUE
pKfFNqz7y5P64jGa/ZGcgyboQGElksDxfxUwEuQzQyYT6wjQe3GaisFGVpav6V1Z8tKs5iub3jHa
0AY7mhNWuIGx7wdBAOnhSqqZssKCRs8HOUxaYYs0W8NafCsVSMVvcnHVaPlVV97q4gPs1muluQwa
hP1i7hSQdrPtG5pVxyekb7UnXMf0J+YdNRJvOLKx1Q/m2jbVCEuQ/zIGo4kab4yf2Kzn1DjGpbv1
1Ge9gD2jvTakoG3bvTto1luLJut+hG1JYAsUqLr+7OAPNuRrgKMwcoHEqHy9JCG+JpRSWFuDQeYT
g99RQqENoqoh67+BH0lwZ2D1GMMRB5MuKWtBdRnA4i3x+unHb26l2ZUfoKk+BH3QveO+uj244y3R
btaB2FBf0W755HJDLZ1Y8cKhQujo4djcx5LyBJsxsKagkteqc0stkj4oRjZSKBpNK441LTn3xJOh
T8ptEpa4OGHJUCfstxRSKyB+ng7wAxs2C7sK0xOZsfCwBfSxjNSegiCb58mhNIxNa2KC672yPpA/
AvVUNIaOYz5wborlRa1kEjCPolXWEcj5kjg/rJir4B9FqhXjUta6faPq4XTdtLlgVR3cRRmvVnwT
wUQvg5n7EjHJupcBIr+iF40dN0bPPu/klVBVv4PrDc8Ip/YoOsht8eG5O/5KSHLZymD+1XSXMaFH
+0RVNCvO6xWagMc7tPHnzLR1mGq1FX8dOtyCB6VGgHn7vke80hyBCw4A4sZjyYdrXEeYTJBkukYd
Brs4ALQMNjAzYhizQKC6pgbPyovx51jtjd5rYQl/H35GVW05ogpkx6P+4uWHg62SZ9cLv5q6jZWK
t4mwDeTIz4b7y7jZ9RQH17QNJtXpIFJb0q6LgbjiuBfo/EqWIVA4oJPydj7iG/aCDVwkYPLzPmHJ
dF/vWcb6a6EcwmSCE45rXGyp0iyjfEBI3D1gntr5NMdkLBGS0bvx7nmP4EjlVfW5uFHqrmj5RhrS
bSvv+7wuMqmXDKnBX+vC5qiQLj93C/LDLCeNR7ynLB8tlKKKV3PZCUThBq9HnHtyWEb+qtb5AZIU
pzB9sXBs8icF9wikSlXr8MDYIWBI1lhfM3cuJCHI7stPBKvhMWlVm3mXZXiPLg+uT2BOswrSaQvk
uSQyOUfX7rumHI0aNUlXGoxZJcBq0xUa4nORk8WcMdHswn7tF0HjqWgRhPKBv44pJRKVAZm77YqC
CrY3CPSH8Ft19qeTVimGpKDiq/uCVVDqi02KqjfeWHMnAeFKKHgRk2H5wlGZybGwT5g/rNTBVv7k
PXefvTIlsZEwlq4vB+XAJULUcXxGvqxmUTToq0npmAdBEGWZyJ4VD8YBc05/rTQoMrTGNgOtRptV
Ja7piZGdjwK2DvIbdVXkxJiRPLDSxwitVLkzeqxpeEwycrCOXxPwWclK2XG6hz8j20mhet/75PpS
Ho4NXC+GUmjPyN+5w+hO+ES0o5mMvDeChy2yK/k3JeZLhzwUuABip313DzebQgQv0C+l/9oYWs5O
ALMz/Nu3a8FGeTfb0BByAF4PCdHpzvNcjuMXPsfcGsgt/RKfdagK5AWHD7t2WodhuHizUn3AGju7
gP4HEWuEBJS4yqseEeTdqMIReTV55jDoq4mJPoMkFEuUE6COC/aFC+0A/392dl8LubHdcqrBV4wH
IZXP1mEtH8LZteFulmDxq6g5waq+AvwBzytsUx/mo9TzaIhdPmtkIIM6rTUp+MpbRj6oTHipvU7j
hRBCM5K+HTNAqm7TPj+u/HaAEfsb9W+pCamXCASR13/shFZflBIFW6d/tU4khBK5aTxZ+BcQZ5Ht
S/UsZeGT7cf9wyXgn28gp3kyUYUoT//kg0eetoaIUS8Lxhr0KIeZOMy8qLnKQiWjjGEdGnMKsU7U
63qOGDLZSzxtxikd3MMDj6p+P/DTxC/WA25vWifrncYzS3+Is8VXm0TkuXFvxHGsV3rDRWJloKrB
RjfjvH0XT8q3rNfASiUv723uLbu+JhhFjJlJjNxRUkYiTPtCB7eom48tHYc6tcp85UGU1+5QvF8f
eu/pn5l4gXG+I/hMRoWJxU9LTvrnBmN3PRj92p3XQ69/hIU2qFcD76SCBzpQqJTT3aiZ6NtKYZZH
2yYHCainwrw/OJtDrEjPemwT8lvf8PEePeloHdEp953W4xmnKP+GgrTYDXIu3fEfqGz6w81cRor3
0ZB4tA4B8MOwq1Y8tK2aJh/1EcGAcskF1v5HW1ALoJn2I2yV75WctzHTFv5EMq3dtIUTWEpSlL5t
HicYwr8/vmtW9Wv29IEcrmC4Mp2lBVq9XYIpX4DtYan0BVOFAx9jnF5IlstxQJJd7U6oRAPjRZcz
XFOiaDcSsRRLUONkv9WzLHxsnxYc93Ti3E6i9XW3sK5y6AoSSdR0sxDTUQjX/v/iO1xuk+ggVFvg
8engeHEnO/0ag2e8VXSUIWJEInYIbPYpgSdbYWImw65v+mY7t+J/zeVANefN8FEE4SGVTYeYF2Mp
iNFgZCDgs06XYvAf5/kIdd5hvTya+5jTbMX2xC3ZnoTn0cKFRVZ28OO+oCFr93HJlfGOpo5LOKcQ
XkjQ3ls4BAQcj+0uwgQCLcz+r5kMi5mOWYBfmRzl2F6SDugJJvGE+ol+V9NdEDgQJWOvncTdvgft
NoTJ9aRJJGsYrdN7gia8lvuqtoP/igZaQLKepz8YnniChqq7okPx9uViu8b5QDoEfmsCkVekMNvC
AET9MCe98+VCB/aIvgI8NpsTP/ZkAdqTZ8JDuZ5lUmYyqii/W0GgtIIuXS75ocGwyQZPUNxmxTa+
Qd4rNmi510yLNaetvlQufk/mSvHPHPioAkEy7RB/AYQ20TMuFe25MSwZwmObd5QA4npOFgtCY/aT
/yHNk052pSLo+1/zcxyHLMUr2Edo5bgwe3fQU0NsQvmnwCmXPSQYTFaEIhWwR9FJBJe13m5d8ye+
X7kjKttyPknkV+wwM1VyXH8tilqtoLuFsACDSlcZgEsc0nWQw+M1XNietlUTj1YFeFeHsxPG+1bI
nnlF1oVhTx6e++2cKZ8wAIDg7BlaDMAbiTD/2gj2tocT39Uzh3jO29v/szw1RqGD/KblwkPqXwOe
rXrxXcXPX/28oQlmz7VHAkINzfurklru7Mk1DJnIcIhOdOrpFoQD3qP2zcTgzFUsM+mcDmizyh90
770HYfx3MdfwlrRXqCSx7F8rgGHVqoEF/L9ZNFMXDb75kv7x5zNfwZAvR7/XCErXPd1iinMeIWn5
b3uMtsrAibX1MKKR0MKoDCkUGGIRwAnBZ1NjQNX2vJDcn2ixwLpmT4894UPdJHEfaGWqmEUtDx9m
0CrOuiWi11KUsV1ccWj58+g6qTHyELU3NOeqxewT870+GfnMI6aYWfHATejFP4ZS7RNhrl1MN12i
gH0mLAPzsCcmuTUzr55qFkOk+wKGPw58cr5jt8mfLhP/dwoCXpzAVe8r6n9nFFp54WLokF+3D9nM
JdQPjM1WRvMaM46Tk+XT9seYVfKaAej/88EOYtw/TeLfWWflWuSJ5a3aBG5RNWFwaMJpq+8pAank
ReFkErSMN9csC3vXPP86M0XAm3sn9xfP+oEbCBIDWxytOvZlL+T13ihMDEgXr5InRXg82ZmBBlue
YIi3QmktlM2+hovCqFNunMArzmcOtsS+yuviXRTQTikpm35hyBbsNd0YpRGWX9I6BxXXQyelPfcz
fxMSAkJDcZHgS3dZpilo0qQ7a3jAuS7bKbAVH6WdGQFCMFYodruw76GGDMb7K7kc/8N+O+K3orSj
ZKO0rxrJNbDFibr8/PCMgPLCaHNaXIjcLdeBU28kleOejtXprECMDfNHS/L/cGInqz1VeORTeXSp
HA+r52VilTR02G/A+PkGq81Byanniv8Usl5DdP+6z2I36HPEE1Rw86dR12sX0UlfbWOJ+wEToksW
VXDO+XiovRGh2raXjcC4q+z3HxTAID/mZekX3Wp26xfvODHGMotFURYWop048YXsfSTViS4ymV8p
JrWCCSyw9irBUMAtU+wmFS7OR4d081sWaXLDQtsAdpJiiYJDHw9eoUllK71REnK3EgV21zBm8LII
mUD7OPQt22mCWgmqQyPygwn9e2eWe3upMSBbYawwTm1uvNj2eE8DZFDxTbx6zmwwdupE4hsw2gyJ
jvExtidlqDcryo8c7x+jCyfg0qGkINiLhMGW7RA8stB9CF+nL1Q34a5IVflddfEydZXE69xTaOx6
IfnXVETo45LNRkb9pvYy7iwLlq8w3iQpokML06R5C0Su3rS5EeTvMjPV5HM+5jkbuSUMJoCvIx0e
08zo/E8audsTKeWbYKMioXwuVUOcLeGhdOKszr2Ec+zo8xWMbQWZ1+nW4EO5Qh8xpTU2aeSWOmAE
MNWCpqoDiCnGBm2p2+GZgenv9zYKveHxgEpVdwdpffpbY8I7L9BStQkEr9H+600GiABG4ApxmlXA
24tqjCsFGC5U1Qhvdc4I7bwQTzo0mrhGNnPfOIIvx++IO5KCejL5TjCanLs/Yt2K7HscR91SZxxU
RDk1qshKP8LwRRpI+pb69TBgePhIrYR7xAvwhqbFmaYXW19oZ9LVKiuKfLiYmnmqFlGzsDXOnMpK
hnpsCDNGOOcgfu5AcNRS9dNZfp7QDVLR4l8NZQt5XcURqHbL5u27lf6uToFQ2gsTROCdFSioe6AJ
U62qsITG7N48yb4Oi5cHA3AoGJADyU+7ruTvJLXyZswASULaD9/y5tvfWmXYLMMuDeHrd44ZQjlP
1V6tzj/5iHso8K1P8r8qQHjnQz/N1PN7ELRvVWXPpwF46Xul6qLLXaWC7y/IfG3uD8gTK/WthbSU
sjxHEcYyRmyx2QITZy4Ayo6UwVpYI49OzJxZb4YxDxmZDd0F72Ri1gZ6bfev69rIRIPtojgAAtlu
1zBwF2pTYt/astSIix+Odo/r/qQKmgfTRQ/5cSxyzQYpJ0UlAdNhfQmBoOGsk5OgWtdgd7LxB5/j
c4r/m4uQo7AoW95mlX3y0h9EhvWHRXlRsK6U0bk1OBcuoHYfX3Rj6BwN7mXQio8/fF34aro6zxP5
/ljPmAnrTTdzDUgWpy5EjDvuryakM2mdHNMDYJp84WN2ie+E1MrE4y+YR6E7PusA7IqSqo8m0gqV
rJy2304QhnluNjcErUBEiq+bHxPWO9PovLhAJh2B2Oiwh6bdbUIjR1u1kkBEZPoezogxyG3D42F2
O6778cfMcOdZRUbfjkGzIVZ3onTUN7kM2jtyt1ih6xXOlVcoLtgrtJBGpjNGhbntzNat8RC7vIEd
5XpBY5Gw6EsGMC0TK4J9aZcpS8ocGFqry8leNrmd9gp8AVLmzVz/1niqqLR1wPOn9OBwDkMgJFFG
ObmXArY5269+BbuMHcwiP/NQZkSeR3Qth5IXY0FJsUnIP+BBbanq5nSV67ASuWcziRonM2fJSXNc
LTHYeHwW0O5psLl9mBiHTu1OzuOoB6LHhcaNm/16VPOO3vT/nJTwUsAncKZngMufTpOyWUhbYxCG
kBCoFVCi+XP//7mTUIYHOf18bJsolEXiES+QCSNQ2SBBj91UuT6gwSdI+1OGGS78qDQwTt6qYy7D
tjLPDssFDrdRJtfs445PSmqclpbw7bKzXVUQrzMZ6CMgZOu7Ty6rTXE0j1GCYrEF+3kHAla9zLwl
pduxel8K2AWxkBRH7u5BNd5ZqM7sXsIn7wmIfv91y1urSZ7l9PvToRnUTm9yblvfQOA6lyesp+cv
IHou36Ts+Zzh8oZmTMcfCI0Yz7D9GmkTnihOM+DpEsqRoqF6YHun8xrpFgAzJnXqVKZ/VL3qFdZe
7dCYp94/wZGcGFp8vcMTLsfBcbOH10Uczx8RGtXKZ1FgElhQU4XMavrP9cpH1ECA+QJF76hs+7db
gscgStZXAQRv2zYN5X/jU8hbAFmOP2eaHp3po77OkRHb6r5bTPMKpVamcUXmGXv/IrzRAe51gFP4
hdNaRifuyUirZkutL61dZfD4MDdgGUbVS+Nz+5toSE7gx6aCWNoyWh2gN0ke3Iyy/udzzpzvNFXS
usVO30BikAjboy+CquQ4fvbEj/pHNpM7Kri2V9R6diFqYyqkPZig+VCGt41blHauAUEzWr2pZK8H
y2b4QEf4Fym3EZMUhzjANkYEV6v+cbvP8gt7xkC8pV5Pv9pr1Ga8Lv27in/RYNv3S2X3j0UgcKJn
If0iUaOZzgLkA8SMfgDUS1aSAKVvKNLDoz6JSNhRX9UUVaf4lCjZAStLDfWpo2dUPbG1lvSCYYwY
sBGMh4cWKfpuzV4ZNcAhvVm7NTuxwAAjG4tYN7KlBicF2wfKtwMIgVF75KQtQ7hoW+ueXyHRF6d/
p6k3zGYKI8pdEJrgEPslyuHwundRAKtobwTmKSVxjAHbkkQxO5iXwtRUEP5qoF/akGAN5mRVomgr
RwnQvf1j4fwNy3oaieL/xGvZnD0a0Ujy0CQ5YL7yfjGKCXakdpj8SP63t+8YYX1i7fxlvdLEv4UP
Ktma7k1wKUJbp2heEMfyG/3C5eFbJmEDo05rfk4ItDgDJaXUSJwyL3x4kJ5XcOYSPYlPGmXt9dip
+sfqDm4xV3wrLzHeqUEpB2gROSL1ZhSLpmUkA/DCaOl9bO4lGPnf//qLi51kYvTFCD8iAcWPKTOE
2kUcRrh8EVWtw/Q6D3Dlow5E5MCu+ZnOBjhfwPofPNYV3SsEx3ImjRslwzxA5a/Lw2/QYCdTKqVW
GoVfVqDMAv/j16+pGMBI2AReWOla0sNuO3ymvEFEdmq/MjE/kfBfxI+S24dIlGVSkpK3oc1/lApW
qgyd6HXq6/p7Htgf8xna2NhAN/KghxLc142XEhsL5lOCxZ95k+zBKBEiiXFq2YvrJ7qplDPkQxNG
jx/9wFvEiPLjVipNuLhA3hcb+AZ0Bdc4nZ7y9p3ieLMqcJfiiMWXSD2od1fLLiE4SAibtQGMcgJ5
qxt5NCHOoT5JjeTZB4Ys86Zji1uX1z7d5mmtiD+Qy4RRd5Q/Q9hhI1U56etbz3JvfI1S93pUrPjc
yPm5YhyFsjkaQu6hGhhn2khnK6n7uujSTMNV7x+3fbla2E7qNQIGd8cBi0YX10KfVrq0+jH/xay3
FZcTqXFTU3CtdVJm9q1rxwjyEsHm4lSspFEwo62KWqbxK9HxAnKCsR9Mk35RXYdQK7CW0/gs52WL
Gq5zzcxnLnyDrSZZirM3/xyOazu/Is5HeUCYkxy9t0sSHBYS4KLz7KvX9SYQ1PzyyUwIzduKKfLR
Dmpqe3S0gl9tjargYsixBI/R1eS1gYwh+eIjMubVqPvapMTLIfmZV3s2zWTn1GWSJqp3o11F0lSO
QrQCn17O7W0wxwU+Kh7UGjB/1iok4BUGztF9i6f2ZNyPycMVOjS3OSXNq5Pt24kFi4S9c2KKXZPz
hEfIdrFxub2Z19BOZ9Hr+mN6CaIx77QAk2RXAhNgNy8xhPNjQfv/1P7uwf+2VY2FjkIAK1Lay+4J
3nTztPrR9taInW5dl9dLek4hMyEi12MiLKRDCyRj3vNHhxKdvbWs+G1o5tKkzySprUmZJagG7Ya4
ZCH6Kv7+rcy/5kNI1Kt3gAvFNwd3rBdGCG4ZAzLgE1DHIGQ2C/0G1BZmJWa69uu92d/MBCc+oJM8
trovs5GzwuN4w9f/oqeC0VOchiAU0E6Cu09ZrKsQ2Le4v/A5Js7aj9TzLbf2qDBAHYvke8KOX8TD
ULEBOxRHFJ1Qb9FgpX3pZb/Zm+ZlJHyhQ5ZAn5ODKhAVjPpcuuc4ppl4bkpMAmJGBSb84Bccmj97
U4Enl7G+K7o0+Bi/LqYXJ/kmICZhkYPx4WWK1cnlYOkTTnRd3iW+dGSVrtVuMGU4BBfCRz5ceft5
7PEM2MmGoRniH3mBhlV8/gMbrTlTrHSuYvciUUMHfDFivyFAnV+UTxudNQQJGQ6jrWlVGY19H2sc
vv6O31znn5wAgkycCTq27n44eIuXO9Gk21ETBIyiisZwhL5Sr4BA6HehgqU8KwYXngdmWdnPlfdm
M12XPXiJKh4Ho7A1zSWb2wPEpBIPkOnLKhzf08BsLJZQuWzLnOUAhf50SJhmn40ZrM7Hyi6UxkbS
BL+eyR3h3RPw2maj2xh2Xg3uBWMFvFBqlipMiq+W1ShsZBFqlq0LSL8d1s+AyoqMC9uj+ttQmDM0
p2FxYArC37IP1/6hMfvHr+LdUJXi3sT1Qm6n2uTfppi+J1WHLkYSwZHmvQBuc+q+Zw95fDDv8dLh
KEzcsD/w3MhzWLw1C6JfRsJN9Uqktmc2CMJjy4s9OIi7rOqMfmd6KqjD0NbgjCssjgtGiIkFp5d4
NMtKCx3RU+0jTm6sysdPyd+eWIMLlQMObi2Ky3tuuiAXBus471bgtMP9jfUZvZH51bpp/NaOIJPm
6cUlXtun0Z1b6C98LmfpMk9xJm23hA3fQSpD0hgDAPOUJJWv8ODzia1etVPuaLDWzpjdhPzyoKm2
axO+2SJ3l9AbqZ7Objdp0jfXdTRj3hZrlTcibnx/x7jj1vhd58rJ1139tMuJ1Ykqbut823Vu8meK
x7VBuOE219TyGjxpjgfOFQQ1sx1aaTNtSM9t2nAESSx4u7vJhpZQW7zT64YPVcS/r24jHjse0TBk
RV50W+bs2zVkUaUsEIc+RRKTTpSlsPkdUoDewBL+PUQyyov6BN3F2V2XlTOOEPR96f7oVqct4AJX
YGgr4+Ew9kpoM4HYz3RIZALh2sQarKhNnmXmJVg91Txu5qqwjL9rDvc4gcK0L7TdXkw9ONF6vE2Q
A2ss86/FKgPS2ZyyPcv/kkYfTRAkI9zjmkjhQKmN3RdIWaXtfqukee46Kgo3q3qHh+3X7LA4dGUR
t4oD5HrcNiSXRM8bBe9KiFulDNxDe+o9dfJ010lmsfaYk3xmf3MRkWHtGU9neHV+sJJiXqbdhfRL
ZNuQsIdMw6J/KVacntx2a1mqVweRQq5Fqj1PuVIn+O/J/0YndERrV69flbys5pK6jyXYuUgwEhtB
TOYqeZFoZne32PehEXpQT4Yu5A6bGXIkWLx2fu+zaEr3wKhSyJYxH4VHp1cojLR5GXpdR6d916/l
WWFwcoP/IDNd7rX9I3FRxatHRgjIEb/AvBH6AXanWH5B86DwPxkUi9HEx3cYe6Nkow1o9QFmxECG
nlSAzz5kDAALMewqX+CpCRfrk3YBzUxkxeDMQVx849LRCkl/7fSy7c7R7iTmGZ+XZP5lprV7pt05
V/EcuUPj+lc+Ud0xP57aRzysNV4VLjwrQQs7WpJdFN3fYfXh6pSsVElgc6ir1GfUfeepIwxmotWz
9YE1LAAawgtB/dFPkNiBwHbXS91ppWrEyB5tgXpSkVg2z5BDFxCT3R6S37VLOAxj469NrlEVdRha
JwscCUBwyc4KDvNGgwiW/3Wwn94g+xc5hBDvxN5xIcyJFzMGS/LjdfMh51HFAO/wSCrE1AqwLsJu
R80Pkbalac2Db/uzt6U6mdLph2dp1ElD9ugH436VjLzYAYJ3uZgDaeNTOQPvf7OnYstykAlLQwKD
WS95I1caqhcdoIoIu7Q6TDsm+bBkZsvMfn6DyZ33T3AM602yTFQ/ywp+OeehjMPJDuSspgM4iINi
FyYz5FCCMJ4nRuxztfYAL7r7hb64Wgvta5LSwveiycXH98k82v27x4TWt2m0trwty09bWlXWma/L
JydM9kxV5HjiTbH8BSbjIjWaxIdOM5oNkEc4JCtQLBDemr3aoTuAGZRtzskBCE+Ox4H4tUE995Mf
X0gBIfasgEWQNNPy7NKBsp570SXmqkQWYTkOEekv5cVVrhnx49LrwHUdqqxiotf5Zdh7Oav1qODE
Pr/kl1YAvN7iEmKgC/zqIcVmGnJf2fn6Gle8Mu1wnnBtiNJ2GeNGOKZxDQfsSV2HVch9dj4Syvkr
cGcqk+bZ8oX2qWldRzEquN+L1RT6DP2DPVzGyoyqNK7oRkyoY24ZJzyrp0Uw3MZH15RHlDHi3pg/
EHQn4dujUOfsTdHx2DVj2KUUV9aePeKafeQW2e5rTrk0NCMSZX3pkLLBusPHQd5WMZ+FnV1gOIge
uU32ZtaynY1uF5o58uvheZymNwZGdPs4jbekc4HTzKodx/VmjX7WXP9hTcHZDj1dQ6AwmeunsaFa
5zsIVkXkn4gUIvFc/7kvlk4KYeMGexn8BWGf08GOO0IBiyCx0zjxSFK/qrDZEAkT9oae1BRe11vA
GlPKPJIrGjhCmm85zlKPNzwxGNWwufL0n5xqgLgFhminXXW2XxZUxKWG9ClTIVUjaI++7+QuqZNp
dQzfcm0ux6OUjH/zL70yIWvBKkcuBb+IEjje8lJotg/gm4URMuKneKJd0ZVGKoE97FL5EY7LB2bo
ImtroF0I2JGOohvuCeTGpPDRKfKupTNoxisrgD2lCnap9QT2cOdX3YqV+yLZ3Lqf5pNNltnJS/Jw
3iGBXIlvpT+vDm2fzdMr8iaJasY9b24syCoh27E9HE7/f6VAs/8Q77jyyi4YR6GGZb9FBoMVy0T8
XD2gS2Sl3fnS132r+021Q/SAvZdEmNoPVwcMbjOii9JU2xf44mp40Ceftiye9xjbOZYjvHPvejBR
3wQR9IT1esw9qeDDVKJRKCT2TyXAUPJctWasQMHMtnHguL4H7c+iGhyMf0ggx5hktverMSjaQBqY
8VLM3LCe0nKF4XNNm/IPjb8TcO1JzuK3DCQGEKST86pCiCQuxUyQU+d7yDdcyK+aSLWi1PVQP+ig
vBHvv36Tqd2uwnOazWQ68Itf07ELBBFMvy9exdPl2cC/NtWp6JKCBRK4WDaHSujD0m41/UrTNBBI
9GIoSCwMm7WDG/BR2CVo6DS4NUYEla4fZiGlVQfptgsd8hxgK5Jh8gPgxKjWmhf249FTCBs8iNM+
O2WLSdXZPfgfb3nhxRhUbv0FWdTGS30NpXeDF3z4B3m1bWR72TnMFRVjU5P5uoqBvItuykV/TvO6
m1sgoZ9j4XsXxO94gQD2xfv5HlJswSbjERohdzKl5Dn3nR/WbwdT06sU2PFVnAy4DtcGPdeZpcLx
Dknu/QdgbI8xPtDi2bM4YwqWWerDMgqeD2wRIDmHRYpY7o+3duEzlOsQrR6XuZ/F2IHwWcvfJ4l0
HiSH3lp8tXN0iyitwYfDMyYvrYzOesG7oQmEFoO6jIcDtzQvm/ENqjyQiQhiZmiWWXJ8GTV+Vw9i
6dllEicKa8wJ+oXH30wvnlG0RLWAB3fUDkjwRP8SQk413tGMSjWp4VzimgvPJb8HFfeOjozjUn2K
wJo2SAniOa9gvEZgp2MEggz24QYYJ9Dji2XqQvDOXzs1cNuwmTiO7b8jrE7iDzrWm0thkrdQDwGc
ttwyak/4BqB/TU5l9SI3iOCNaK7mDQ19QiCO4IF++AqOOOcG42rQTdUp5kslU0O0EgXp/qE5g59H
j9nPvvJBXzkohkViuSTU7zBX6qH5mJ9zah3uduJCN6BpMaRNb+wevhFzQdtf/UCOmNNJWhr+72zX
VH/bqcJHBE9fTXQE7SjzQSs7uYNUwfkyEGu8FKetIaW8M5cZeKsRfllTD8o21YumrlKizaqBb3De
JxfgfCWR23F3HZEmIM+jRa1zwr17kD4+v6bVvBJb7LIA66esDdiyIg/d8V0cVi8aQBLqMfGnfxyg
TrhOpj252xEx0gRKMWBrDfbpE75xVgHUTE5RRnV1aKsXlpkXltgbmDua/xRHpAnJKpUpacm3wKmY
WgkgNQ/r6WW6VTRO7fnpK/cPRW92YFAGMHQt8/HG9mjUxA7GSexEgzg+UUMgqslCAp6VOCcVO27K
/JqTq7jLe/QJnechJ6/dTtuvn8UN/pOKxpWOCEhWzki577CU3F4t6G3gywEeszkbOmBDRGCG7z79
UqnWpriA6b563tH1U3wqZqqEYIZYzXnDSOwMg2mY1kwnXoqPi9jteMmDhHl+eFETUiBnon0mEGQV
49J7T5EmIdNR40QGqbhcl9+ZvFf6oISMjfIDubC08SNeV0baUw9XR5RVCZZyaRcu+qI4qvNbTd7T
M0IOux918KwNsqgpx+urNfGCJucSyt3lpzkb40mi8FU9OWPwxpMyDOgt3oQyUa8bhh+Y1UqlrEG9
8/u3xFp7LIQ5JE36aauIaHwI79HoVopmLqDYQFyDXmxIdaDxVfqs6db/fDxhuaYZYLwm1Rj4ycu/
YdeHONwQs0goSB7oTy+cY8qtDAhgvyzrzsL7WWTIPq+OqX2say7BxMUf3v1ASLm7eXd8Xt0baAxl
k1AmikxCRDqhBf+H2pIm3/3K0TlDens+UbANS5J6SXiKNyyRpzaoifqlI5BddjhuDdczf7r4i0mW
8/IVzYL5K3eD9Yxy7GEr3a6jRmCIujAUfNUhteQ5w6MEh6tv5hoNfDTU2ykiIZJ6GdamrazgkjUP
9dioBZA9ylpiq2MHMATH7s6Z5Nmf36ppZD0dX22kfIsfcIOW0CytHT5pFDnhD24IGuscDEkSxVuC
62cMjKnFSdpdTR4pOjgdVHAsSLcCAXeCON5TtzVZOKI5hECnLkTii+EBJNyBN52CvADgIJPfU+32
/RMQYSbmUyDot9OsXP1tT6HFjYWjoqRe/B/BUvZgnP41Q66mnQdHQwMTzvSedPLIsC/TweaoPbUd
d7AUmh7NKAAWPnFxDqVwvwIuQ3B8f6h7Rvd9KdVv2ZgxgWvwcvsztunFCQBGwwbI1+dYPccPqvpa
GUUZqYPQ3KNdTlOiAHRrSAaU7TQTGOEN5reJAYvEJW8qQeOoD3PoU6x59/a9z1PozJxSCAgwXwFz
vgztxmYGQkcdMgxoPdB74p8G/KYjQDwGlw2MKlB8A+0Jv2Mzjs9GJzHqZgUWOzHnJ8IDfcPjf3JE
kcoHd059QzVgW6NSu77ggP/rNMuaFD3VGZrXxv57Km6Mi1BbZhTa5/bAXXlGxf6IBNFJBLmM4pAZ
QMgdjh9fHsjayz61vE1O2Dlvp8jT15CWs0hB2XHewXAtuJxkWRM7kuHdnPIA/TFlw6hStZXcoX8x
epH21oEuaScCcb7WTz35PDZoKhMpf2JyMYiCX23kPTvQyGNsFsOotoYP9OLehnbJv8g8i+WEJBhk
6OyVRGxQ1VKkM676Sgb+g0uHNnVGTIMbfeXjx8AiJyb1Pm4HFJw2wD16ghpc47v4rLIyFC4EEln3
8lsyZxDchVLXwBVoRFOJuW3ayfJmlXIoTX8NXgOHZJ1ZoXxEB9eagzNDJcWYVnvodWqvywfnwGyh
4/x3xm22epMGu9bHfU6ra7aj8i5d87JjDR5K/7RQnieHjD9qs60C426SyCq5Br9w3tFquBX2irlN
j/oV2+WANgaIarXTzNujgL/Fsbnl0/w4QNPraGx3nPUSwfm766zqj99w83J2Ks7GqN8z1C9WuJ8+
GbnypTQ7iz5bAEMRzW7wcieNIvQB4jNboaPYe5PzbMlh0aticEHDkKUYqvH1FgkqdGXtmNGUdkM6
2bIEAEE9ag6FBluZ7rRThILVeliOCcQWYkMWqaS6vRMfLARuqw5uQGWqZeOcA4rstStsdoRPxpu+
75NCSboCQos5GK/1iBvvGlhpYYnycex9YW+HSTpBGk4FtAS5EibB7P37X5IK+lseA21b3N2UX0hM
VSt3Z5iKIm83Mtu0wh2NYq9nr4y6kJ/Q4GKXD+6d/G3npkijzhdX8s9kEUN3bucLS97pLscKM8T3
zByDYzV4OFCCOsRppTt/jpMi5UZrRk0lGup4OEGH+Ha0/iZAFpwS0Gp36jF0uQBllzewDWhCINgx
89BRUBxv5OQd+JBC7aCYSaApqdhc5HpfDFE7UosDxkHix8IPx8SgWTEC+7FtFLXprXOpVKJ0qd5U
YfS39SiHB5aLfmjsHDr13BLFVyj/zjBvNr9okmPZn7vhUZBPs/lQv7crl31R7v+SMYrfd2V5kVSJ
pTxB0QirXT8ohFEuklOaloLFltTnEVrIipBw1Om/yWDLesRAZllXY9XWHH6wwaOwl5ar/6Myj1UZ
NHdtGVadCcUGShISKdkQZYE37BswoDs0lAJSXjll+tZpFypfkk9KAqmckn8rY/JYRIzhs69ZHxYS
u8oTyjzlidR3FxwwM8Low1XGs8cYtaEthep0lbtiuKranIutp/ylrpoXKnW8jBkKuyBGWD3l+7g7
HWI3bst2ega1EHVUfMK3By66GmMpYkt53Nf0o4g5gqXynOPFxu/az7cPN5FXdBWj4o3uhpZiaI1N
k0iELjn+5zfvsaAIvyGu58I/q8PounBHicKd2jP0NpFKuh9pAjJNb0XAW1zhsj9tp9KNg0H1z6kU
GlNtRVyUo8WG0x9e8UKEU9TjED7XbyAm5wQXq83pCOSMZV/15l1wdArWWbruMSbQCMw/kjOXdfv3
fhkvr1krp0kw1lxK8ikonMjJn1AYcapKd6XPYM/OfVjHiIA9uvM8XscFCSy7IHfjetPVXGvUv8IC
6QHGttvQZXrYCMERwY7y5FjwJ+h5Z/UTvf1AgCm+i6FIsxG+dMNfldCH+XkVeecUSBUsf6IZaQ1b
9qOhvlJFpxXaQouWKdEWY0rIGlumuYHCLk7oFmkWv6z75yBLDkuaS9DgR4qIpOS1fYRd/5/FUv4c
5mN1m26VHQfWASe8SwFMx/2gwYG6QtL108cNeIqSdex6P1aJbJPPxmJ1SD11mL+OoSj/yJ56KIE+
Hd8zXbQtyAWoALuKcxyPKx6hREjadxQohPiRhdflrXVjzmxEVo7+dWDy5ijc1nJIqD5rj++OFk6j
DXpP1EPppWmbu2cNoyx7cGSMwE4LmK835Ea170BVkbJoqo/gyzcVkE5myQxgytTwY2pNcj3LkdHQ
P9B4gKGoe6kFEw0/3NuGaOR7KKzVVPhBtmzIRsYC9Xsz5oV4ygTfRChsyOWAU8ev34GQywUohjtP
8FsA3Qfzpd12nZ0TnxqDGQaY+xXJ7nIOnN8D0NsN2TqIf+4vXCgzlOoYkeSMHuia5d5aDKTSCaaC
fmbr4IV2YnfknEjUHHRpexs9HG7cYyPnTvGuZBdBmH5ogFIx7mN4QdRJYh56lkdn8nbe6X7AKas8
A0m1JU77kSClHaBAYs/IJg6l4Fv7OleUc0hkZYM3yA+GiB5Hq1syMN60Y/2gSZsivbmfQ8YLXd3U
Z9q8UQ17I3L0AbZukkmB+sjZ0LkiSGY1KXIgd+jQ9Z9i9TD8uHBE+fGDxK7uNbWdeuuhnczlamCF
9YJCp0HPu4RtFlQK7DkVf/ti68XwTPEnVIie/AxsBCRSHM1e9NzfTR6A55bHgAjk/yf5St7ty/1W
2aOTdVZtt5mrhAAeNEhC62yx1zjkNnVX6ar9oG0p7HYQus8pK9pruZY51ucLR+d7eDAHSL+FIwTP
wTmYQKrK1ZdOsiEv4ad66asasNBRT8AXWNvx97NEmeB9DV6rAUtFBhvRAUE94a8kRKujKkCZjwO7
p0VjDogW1Y1xo8PKcDLsESDJbpwKkkw0bwhg3kyO4m9+29jI0Sj9KJt+qz3FIdKwhP3kRyCWpfbI
LEaEf9r/ry06D7RUQhQqF7fTTsxjxNSYMV9k1uPHBX+JTaPvHjjJWv2kiymp0O8HtdGF3exM0I43
AgUHZnuksfE2b1xLF+6jasc8GuPe7bb0QoaYlqM0LOJ+PJYtXblz3grZIVNSkCmheUOSpZk1/gdV
c+fcWgM84N3KS9xpkVclhVpMFltoK39Pb0YcHHVWGvITaQNXAhf548a8Yn/vHp0SsQuQCxtQ9bGT
x4F+VfeHkazgEU/jP6DQwkaJxN6vaLDOUp0PK7hGZLnOjSyXDmnP74ItG+e7XLGemt9GXsEpmsVg
69fuQIpAlDTOM642/xbkYJFiaMIbwmFHYZMCx3SF87YDGpFuwmBoW87IABez0QCmvdS7hqo1Tcmp
NqkNmwhV6IVaJuulp6wv8zBHQG0HNSzSoDB8lF50TC3oQC1zq6NNqYQEKe94DOcQwFpofHkn9XSD
bJS5PWWiN0OzTfm+HhDzs0L64M0hUgyL4Z0NZiI1ygg8F1c3O92zmRKPKQU3qqRgqlx3qETd26Vc
aJF9ZCswMRzlrkXMy8j1jxA0T1+j/gubiAGS9dfHWlUAMP9I0v+huccSeiJNnlf8mX3vmMX799fW
jqJk3tDckQ+e4r0vJxnZgWSwbTbpwo84mNBG6A/5RNVH4DT3dr5gt7T9OJKFQKzftuHc6TAGiDct
SqyBkueYsyfcJB/VSOMCdai5ef3zsPeAO/qkqVUEvA5QUENL2gS7II899KeffqrbHgZ9UozPiyl9
qDiWm05QKs0H3TmTujxc9j6d/8NWuIBCGicrBUXpKtocjvzQ9+cwNDkaF4xqeKksOIqR15di25xp
N0xgP8J256qmDwLz/Dvr0zGsB6FiN1VbVAi2CPRLn16XrjYISJghMhi+bAIyIxJ9Zb/COsjIGk2D
Jlcdp4bU++5VPISmmu9gFGnEEaauPl7ZwwJeUv5w6p0A4/ghYoaRiozC7UqyM2cy45veL9ardUZU
cgzaCeIGsFVek/dHG4/kfevkdxE5XySe0CsP8YQ5kkzl3gy1mfxPWAKnB6JSTZ8jzwi6G87xBJJC
tfCn1vGE+U5mrLz9S7TYWEFbrgqfT3D+LD1RN3RqIAqUkdZvc+ZvvlJzDCuiGUOrfT4ul2eJvboC
tEWP0u2vzrZW5KIQWxJtLikGLcYZdzK0kjTyZYJHOeY7LFmJv2/5LuHh+iKTpLR7jtUH0wGTE3LT
qUnwVAgGiv2SuiIBDQWjcZfARN/gLOE05y+5FCSGUCxc6udDFEA9uGzM3GNG0V7SIa9yT2xkOW/9
uyNJcuzf1itA0pQFwZF9nbZrKrKpw0AsYsHOxvayhnI7+riMuEsXLN4e5XG+jTXYWlAEvDb6TlpB
JxNeAejRlSYdLOTjR3z8XysFFOUeWxdS1e/Ls98mtHuXRmfYyl4ntdv2EjFU/bfv9rzhBKmtKdtj
FSbxMbbe4UIpG90vZ9pPOPFxfX6DW7Q+g8SxJPuvZUjvQjfBELni0sftCY1C7cB3sd/OZYgHXjwo
4pJtuhUcaflCAzAWUbHP9OVTmdWVHZChC5ovuVrHCFVYJRaUOIG7hZy0FLO22uZrpEoApXk1suph
BRUKL+la7OsogQ2CZhRtgEoush+zK52D4wTZd+HJ41Cy5s8YzM3eox5/Anu2LpieHh1syBrvvUsd
/KXdJSsS+hOlZSLfJGtvqs7ysdsQSTrJm+cAfcLsZ7p8D1Pz3ue6H+HcXo/PzcukwAnpn/bHjQ3x
0Y/IVZhzkIml5WP4SItqfWXyaoqGtQ9nA0Tp+7ZvgOwKANz1QoaBTfEpQSWtaNquEtslQ0/KA2FS
CjmYQBHqPvPh8fh8A0BHNWMfmWuwUBKM5wO2ogDmibxAtygEenpe+hDOv3bBvn/c+cun/GlpO+kB
UnM0sL61e11n5NNKJpr7h94CyygcAm4LM4Aspa77zCLpP4JsvIlM97RQCO4ymiccFun/GuLO9JlP
A+eIDPRHjOiYhKhqDgLkg88F7lysljzIDsv8VnGcA384LF6cS7Q5PfXNaRehOu5M5k8T1gXD7Z7d
M34aC+KUgRsghcpa00Ce/SZgBx8s6L2xvK78b0I9ptDX3yPYHSGclAiPpzkoL5zjuclFtkHATpJv
8xm9bBX/dVHH6D1SbG0+wQSIkmpHdLE6uKjVgNaTg363N7GM+BPMC0Xdt6YjhBA+tfEAR+hXRWKY
GROwtwUQ9MQ4BOtS4rydcAFYFSCFVerKABjOi/sl2hJLesC6sL5yPXqERIT8UYK+gpVG5dxfnqsa
CbyHc68Y0g7iBoim9afyJENWPG93d0X1Bbetr/vGdD292AyJ3QN6Cas7FFyPHab7Azsj8MYHhxSU
smJyNAw093PRHqpUJdhacvVRhY4saq+vlwjAsBL3MT1ibtPI8m44wYjezstPAcHU7kt4wjKuZkZR
0RrXIriyfxfEHyBZzg1KxxKaZokSMHlpK0fZ5UWjXLhFLfppDUEb8pgqRlKGHc/wsTzryLf0SqYX
hyZ3/jsBmslO85dKw2TO0CilwtgKBa0uPZUmDmLWA3XPGI7G+zZ8O2rcmwhdPssviy0aqqj0XdoW
SncRgMVe3VphHP27Pzt9K/XFl+pbu/C5KjgQHOA83RxQK8pQSvKuhlnOGQzcH+I34Bi9Szge4D6K
hJzYZR6QZzXp+n/sk1a6unJtnDPHc/SFmYi0X6FWdqOL/cxKk8QsJ3FUHoFpSfjbGlh+/ZSSBvho
JsUGI5kDXP6n0X7w2IYPT+PIMIjoVXdp1TuL8WKP7G5H5gT/RIguhwJiSCGlexQISSTmKhkiS7rn
ddHrcm3tbFgPQa40ERsTwDNNbsQzk0EpDu5xOH03ZIkDjOhci5CTBFYRrf8khBVMMHwBMIy5l/QS
LB4dvFEco5i1f/IVkNG6kN7G9OV6X/r7Q1T4GMZEnqz27xZhErO/Nhoi745CE0u2ZKzMTYteRFXA
/VnvotJ5MfCHCx2YQoCn1ZPWLEmJrk2+4AehEDMbRhCOvdnTiqMMq7uGm5jk5hCrMokfvjcsKZF7
254QIjVj3PGZPIZwUTocpJI9u9oMKQJYew2/hqFdWxJYvau5dyolwm8luwOyYBU/IIVAzsoa45X5
yjNOLkZBoUaYlqYZjm+VDF/GEZ/xgu/a7388IoABcVkFpK2T/WmQuDJApSxSoOqwKU04e6vA8eoe
CPbY6EfdzNJ1j53Hp6qF3BbGbgq/CeLSLiJRd8a0u7JTn5VBem40c7SXAttxJ7p0ONGKDlgkd7XP
CNKtYcbSVrtlqx/Y5RecKd4Ye2LymrCwpVHI9n2dM3T9cjRGjYGX1byovoH87WTBdcnGlPIVO6G/
z3WLM7y77banHv1knT7m7AAvyMZm6VE9zq41Y8hipnI+kMGLP4U3/VxCXCV6xIf+mZFKbX0w3kf+
IVYMDIRZVhOb0LPYpRlioJaHfWKwkeRABkgaSZpf2tI4QJLhlGwFWaat+Gebx0lcYlVL2B5CX1hA
b7j8olwxlWsfk1dBNFT6f5Vef1dGP/G/ciLDZWlcSvcWB/Rkf4gS68wEWSfd6o9Tn3dtSZnjSj0h
zRAw9p79ZJOJ7BTRszgCCQA14opIFAGcw858+h8a2t8fm6YcC/XlRmL6L3kV/GMn7Ud0M1YTc0V4
QuuCA+URQADmUh0n4OcLRU9j5RcsPiuA8Z9xdh0sfR2tn/3KMK6f6pF7kArTQ66XZBgXf87HZO3m
4LUrSmGHrc4a9NLqCPUtE3OLvfUImUhYqYgTmFdkJ6PB8JsoR12hTCCOtiJFCYLqUBmZ6TRDDbC0
tnVtgWOV8/vP4p8cfUJ0u5WLabg/gtHYbXc/hF8OAQOX2RvgdlqxxuYQ4YkQpTxn1CFDxndmS6uB
en/FyT48ZwP4M7xvf4RHdz4Ky+0PCNRqycODQXFztrwdNiWCwbUbwYwV6grQ+gztQUOeXwar+uYP
Ux9kWBtsJJ74KBpXW7i4PUadtd8FvSEvBuu/IMXSIk7I9wIQnAS1KVEPjZallMKVkKukcjiUpq7D
eBZLwReI+mTfLU2szPtJTtKZ2KzglSP0brB2GOOeJDXTY6c3skCmDTqkwvQ9WgnMQ6lq+cAWW5h6
HH6USsufXAuiITnoWMNvf+3XAWO0moICuZ3GctrhrDWFz1GDOLnV4clCvXhRQwz/H6M2bR0PuWsf
PzPhucB12rjurfDXx3gLGP+n/pOiMmm1W0RE5QJrvLV8+kzsp4fwAa8S+RRQVpi8lW1+WM1J54Xs
1elVBA7ew+q1gJkJHWC9vNiIHNyn+/abLoTM2/+9gtxS/xblHp4IN7dzblOTa59J6cEapL760bGe
eZKiKX1szEfPhAaZxgjanp3G1ajLKZhgZ7a/fCdIazd6EixcHrLe3EI//CPDFMoXmL98HuklfJ5n
Zj2+tdItIrJyjnlDe5bCqdT3cu0KWOpWOdD1zlwuG+Bnm5Ky4RfnMxu56JvNOaP8k/GJiDLw18jt
uax8DxXHrweGsCWt3rOG2gUPxHJxZ8dv+DdHzTTU4ciI6rXxdKcIf/gUnD4Il0VV0pR27puWVkeH
AAk4o8CdahjL5SdVks+wEY2nrnNlkmnizZ37A6iRqRRkT+hkj9CQkz4yil9dJtwTNaGle3f50Hud
4w7Nk4ZzFFcMIMsyId243+uW8raw4hmLjv1nZVVkoteURsfLZ1H0SKdZdvxaR925VsoCuzb0FXVC
KCZdqzjJVeIhQxy9OxOrzunBFfuckZA/Q3zKsYWgubQk7Z6lsVV4OCPoAuhs5B5QGoL8u1V8eJ1X
Ge/k+JBWmmHCr9xDEz99fIBkBA6nODYvTTorFm2roEU6ADBZs8ZUrTzmZcrGG/C70eYhikodPI+d
jbXiW+6rIv6doDD85Aye1e6YCxSKLxCxMoBCuF3Kdcy3NtpGNEmbrLXPb0hWxZ/AzieFtTJdxvCl
14FJqRR2g5H8pbcllwO1p4mHHuARxX3NAWW7wnD+1Ln9yAuPvqzj4vFd0BBrsa38KQxOEhNGI9j2
IoM/zRNk7t+xCiC9976kBR2lBmfjLYuOsRTI15xlSYrBdEgfnsKF/CJNtslitOVLq/7+M5SG/3kE
dPpaSWvQia9SyQnXthd2UFmEjBfzQL/hwULn0D+Nx0Ig7kvFDz8UN/JS8EOU0oyu1NibUU/0uOsf
5BdREnfBNzFU8XybtHHt6DVH0JZb/xcdc/bkVS7io6K0buJVakyxMstS7/HqCCfdRdrxbmb7n9wt
yYEmNzfGapKl5GVaD7HEXbHUEKc3pQsTgLr2FRi4UOfHmVtha4k62soKoUTEcDE8J71qxb1+bzIU
0fT1ztrKDshK8KCE0/WZnZnx7URRPm8/No/e678iDChKZVvUb1xE27w5c3SJYG35/w5jKgd4S8yJ
WrsRAXBK/YMmbJilpfXkwAMO7paJ7eB7ZDBpi4LXTVWMajNqPgcbC6Tg417KmiDSaFLY7/3Twh6K
fJWpz6f+W69HI5gDNPzeMX3kLrwDIL7Cs+6+DlYHaxEBc1LI6C6ghA+Eqf3EewfbDBsTrX3/w1A6
UBfx49xcP4/mWsMZ1mIfgnYiJKZp6+Aez/7pkxp7jVLhEtYFr7JmN/bn6H2JIa/1mp77ZWXdC/NU
UzubMsv3jzhul6zxxY6+hIDsW5f5/pcMCRb3snDDCFeghgLA0URwr6L20p8h5/sutrhmEfwzBUoD
iZ4/iWZDNAzJBF1prag0KzUtjmY7sHMrryZmwdcmhVXZzYyMeXn2pXaW3Y/0ZGLe/vdF1dRIeQ7W
PplySX8aXjWAZf2+9OFwmi+wKMeA/BQv+XkvxRvSbnFDsgLnJp0R4uczyoX8muBJpTegKa6QQA70
FB+iDJUWlVSZbbWQkVzlFhq9xBQvYFio4sEZCcKWg+MWZ6xcG3qfOhLRqiBWEURsHu/efCMC9kMF
f+ZDmqRXl94JtVmhcqiN7dg181/Ps/tq1VVTkZ5McttMFd4gBFl1et1HTJEWVP88bGajZ6Aivqwc
smpDbw2A/k5/k4W+u2QsYHFWxypsVfTbjLqcGyr3ABQWFbd5KRVl5SPbg9BxLb0KKg1CyffnEalC
lyltflol+wtmsd6ZkavCjyNY0gwSTWOxoiGGydmfmCCgFBUD4rTKG5dwcj7pdZf/D7zwJ/VpZvLd
V6bv5BxwunTp6Lj0Sm92VxhbRZ6+XRxUtsGfwZlCXDwfIYa+WbIFXbTLHu1tZdkzxaKLg5SXry1w
yZ7JvKP8IamHB32xo3QoPQUrsVgMkHqvE7kgUCC46tQPGZuu5bWJ7OU/icUN9mkTxtxUv9SAiLhy
Ang3UwpiPre8HSqu34FaoigatSwvdraxNHECdePYE8LK/ZRlXv8wPI/EkGg6jJt2IcdcOxYknLNI
BBR5tmcrH3gcHdxBLA1D2G1om5BxecwZP1EzlLe5WlIWuW63q1bSf72J5PyB0L/55aedQpJUDXaa
a5R9CcQoWBWCXjS32EAtd82YwbIsQvKdae1d8/vZOLzfmEF2QDtikCQWR2rKRmwGBsMeOx4YdVo4
j8whGuyBX3tRrI2qmyQd6Fzi7ntZP+P/ZgkymsBFZeo4OaMuMO0dhsFt8Q90GMDPaFZ4DIaIywDp
jyFttdlQzw6GZZI5Qc/Wrp3PAtf5zjRxyhCb7g7gmPBqxDNTolABTCw5yQkMVZKIJaT5g5dmPnWz
J9VQXhUlDhlG+v2+7Qpqi7nicZ3pg6N6Qm05hq0M4c+DJPM4/SZEkPXnKzSmJYS6tRfNf1uI7+to
b9Uge/bhQYP58AwYpRtsrzFcwPzMTQiADbVUo1/SrkRmz2v0habaa57aHfdBB0nHRp0zkTU7wkMZ
S5/hLZzjn+B5OEq2mwISxZaoTkKSngIO3S01/622XKlI2srvdtfv9NtVMQGoLXBGhQkZ6x8cEQS6
jljXLzcO3In+t/MIYU5tO32xMKqkhXJtFFhCV2T1wNVBr25OEcGtrIqAX4DkbxdticI+nZy+pqMQ
gaPD/r80j1RFlqTQuSHIk1AaVl4WLJNLxyGq5JkwVat3UipfVdVd1Vc22Nqp0FPPkCItXHIKrBp4
6RTDngcAVzgf3Dpp1xdzjs1gw7Gc/atTtCIdIcO0cB1+i+CCfm/DENmV8vCWNChEj13Kmxzxa1E0
zX3r0F1XJ0n+/lfPSwbtD5tKMeN/L+GRw41SbK78GPNKF6hAj++RxkEPS/E9FC0FuGrZzE6Y8K5p
k9vaizgEs2MlwEuteaFyKZRkBZkhn3W0v1OF6yh41PRoPG6oQGq2GU/rLXQ6Kq6tDf/RtjbhC08+
JdtE6lvAr1hIzF9McVX2e+SIJgnEl8tSqZ65mkTUdxpKleRgLjRXKuSg9/AfY3PmX09TDNOIX0k0
31AUU0g6P4wY5BFRqtOd0yL46aaP1Pv5nn2ckIgoEZHP94EGAPah5dbzn0MOZkAYQZCA4AvyDObD
Q8L6avd4tALQURrM69Bc36OiVPWfY/GqA+ce3baPwpGmrg4XgI4Sdra47mIsokq/cA51wbMAXru+
0BfJ4EX55APNAQLOHpW1LR/H7R1fQppdqnSd5rnsCXmZu1zSL2Xw5tq0g/JT0FT4l2iAuS4I4RBI
ImPR7kvgSVWzKeQjSZL7sov30P4BODy/S2N7iKdq/dvHIBVYkTEZ2oR22wBYSqD71hTbn+Wj3nX9
awRcRzcv6O0HpGQvKgZg03TdHjkOktfPuespN+sui3Eshlff11LXRescpRJlnj5YKr5AX1ohBCBB
EaFaL2eGFee89tRVNLOLcEEFKpM5yvASJt2ZlgLedQKM5d90WYp0q76Cy+LU4jN62d0KPYc0tXk8
Oachs0O92DXXwJkemVB6k4nRcq91E6OOVZL7RryVJXsL1Bgk/X11J7eYxpEuz/OFRB2vHe5+OB4k
gwIZFEqyezK4lBJ0jkB+gNWNCSZFinZn7p1uXDSBMGj76vSYGJ7hKqJljNi34zMqJqE8KSk85EiF
C2neHFGvUkZuDt/F9m4df/3UsSKe/KpzELurcnjj8z0VmCKRz79z0dAnONDTSYpcl1O8f0yt/aAc
y0CKdnem3j/zkM6pt/QRUGGLAsIQczq/3XMCdIzNgQ28wmFUkid/IonXeU3GVa/Sxan7/GChNTVF
x5AUKfeZXm2iTIUEfkrvLBEn7P/3yL2Aly3LTmbq0e1FySPp4m9PRbvPhz9rkZUQK1Sao5oweMkc
DkvoD6BPZbrLlqTsIY4WFTulQZWUU9q/9Ug8gVxu3pncd7+pdQHKIxxjSj4i06MMsJuFG+AjbyG5
HZssjEz5ga+JKgajZX0rCir+p3gUuCzPvYKnmOM+MxDu9qJcFMmnhgaVXhdwo3GYriXW05s8RsAK
or7ahAqBttik5M/DIT0HAHT1V3uVOtbUeq2ZJIRpOt/S1CKysfuEwwLUhdo9NHNOOzIeCVUGYBzv
pQiQN4vQ1lUPdKrKvOEZiwYi4y6Pu3OceX+JkVI4YnyeoWHjMvgQCfY2fXCSYPfGn6W6dvQJw+/a
1SCqXKfYDUvA1Mpj4UsRQQUPartQteFUlQ7jPer2gaMSwCX5qDvHI2qMWFDd420cIqY+44Bl5MFI
9i0gQ6EQAzxo46D4jRuZOSouoBfBiXAY2V26E2GTqER3A69Tbf5UF/jI1YFFKeviZ+8pDx3A1dSO
TURNZy6uf7X9R52RZp1auPdVS35cIMSSzXhlmfjikJP/uSzFkA4BS3Ma/lWE44tOdwn+NordnMML
1Y1K2UNuw1HQSwDx69ZnB2ZGnra2dKz/Jh6haINNjft4Smp4gcV8xBmP/OYYzRH+lRm9NucOECNa
0qXeVEKrN7ulbJKhtUv8gKIV7gP6QUIb4DN1qgphcRoCUVbA6gUxVfUT+CrnPRCBEq5vCPv8bsjI
dUQHZlQdkn2jm1/xGACuy4ZGVYOTW+sUJQt8EJyyjTEkmZNWeN8RmjVY4grwuqu4hdci0DNG3/2x
1EuzG6JgK6nd5uz1oehhegEBVwDLq+izEw+x8yXiRwpqv4ZtmYss4Y1QS5B6grEpSsxkE4vve5e4
ERmFHEFfrnHw+eCKJ2nqmv/mpu6FPZpbOovXy5EPdhXy2LnWFZaDBrXTsDuY430xd0j3xQNviB5N
cSoSkaP/Zn5H9P9+nKtyGgUp8saQ+hJ/H5JTIaleAZzIboP2a92AHPLV1sPcbwb8WMoIVMIGn4/L
lafnehEbGnP4meO+WuM+D4VNiPowcIG5zhHurC9VOZvlnU0iLSXkmX2NYfkmTGk6nU2x1FkDBqAK
tzxJpGGNBwTBHWn/I2rt7V7JYyJyhMgNicozN7x9ADdeIoD5PZfl9NNNuhG4+etr+3Keu0SXgQ1s
gl+yuDec89shhsP4Fhrb1YF4+O+gKEL0E4tHkRfiZZib1mEYt9UpzbBLfEXW2L0aoFGYMW62wiVq
zp9H9/0Ng2vV+6Iq34inPSRVUkWSFGJ+QQM+LN7pFlZTbHa8ErfOVNPpJdgDUgz8XtpXCAd7U3zV
ukBcxv5O85p4iL2tczMNa1baUKJqPM6vd47nQy+5vzgofOExm9A68XSyS2Yk6PRUI4Hr2UwrgUi5
Yoy5DU3Bnvgw6vNJPX5SVevJnFOSgTKz+uHem5OYW1Pyb1KmNHZ9V1StwuVD1I/YZgUfDAAozmzl
QjKnogCkh2p0SLx3fGId6Gy2pBjXKV9rrdpdPAttBf5//azPkkpozc2U4FHlwI3x+Fx/0J15pYzv
WeUk1ds/iSx+mTWUMdVWJfabftRTLC2uGobnviBD16IZ32/nW+FnCgLytR9HQrQC19E6KuEAvhsh
/EQgaS0f25392agopiNt4TsNYWXouGDvWYEvltB3wqSVoX7Lq6nu38HQ716/nyuoY8AHnRdq7CzS
MMuPjr5vKSXBZmzFZFM1BTORvNjMsntAi/NFcrH0RVtEQfw0u9Qqjtj+kMtLzxd9Y/N7FGN6DPB9
6191ffFCWm//fi+UeC+e9lFBjzIuKxL+XckHVepwEisQEa38UNHLdbOLS48xMico1SVIDR7YgkuJ
+QRkiNd6Hi1XSfZmHd5vUW0i/bQqdMGiGW0ya7QTfTsi+be8QKD0GFw6APZlDGGSNn3I/k6TeHut
8wjT7vatw15WTwsqyDAhrVmmgN+vTapKb2ASW2++QClBFQxXxh5d/t1HErDS9G6NZTVr9rQwqePV
CciFFmlIFdlQhIuZBbTTueWHR9K8Cp9MP3aDL/vb5Rgbat5hOpxBhTZp8QAP0trUvh3w5Y5yLM/f
RpFKzm06n4qVmZEibmm4TpOur8Vd3hhRmrj7Y0vYbMbB+6gKSZAISIR3xpyXhDeDixbf4KtPTbej
riD+XrZwaTLwRmhwLUEVVL0t2hrjbeRtGhydufuck7BjQ/d875VHOCS3VbVo4z7EhAu6WIDsNj1c
HvqtsxZy8QzxxG+R6MFofmokxDHHpmHkuyT2SWbUY5PBsMyjAfs/2zSM150u0jFOQZEcA0uG0nw3
JRPDAakYx8a46RKvZkvkATGQgUwUFrEFfMoritKhWjborqgJ5Y9QuDBbZtaHLaKqW44p9RFDOUu9
JKGJRq6rhXV+2xtUBNrrQqjBax0zl7EUNkBkZKosv0UHaGMYrWf8bhikybcP7BbDteUifJSpQVp7
K/uYlxelDdS2ObFmd0NcwjUkyRy6PBeo8fsVFUpWae7JQ9VDdp7PJhihBXZUf5JfSn4BiQqveAcX
JNr3vXU7C74XjJLeIc5rGBPAYe+fG1koU5ITdbTSi7E0DYAnjFCb6QZ9qtS2e6vBcekwfV7tYgAW
ItzQcgeMZy8sAP3Dj8w6OlUFk4z/G/Xh7BPm8ppNrzLjptue5RCAASkWnPHLgQ9o4u6J/ynZjMK5
9GDcTVWJEAPou02L0xY4u3nd+AjESHcfvR0nCqD0TBgVURTy/62N4KZM11+AT3xW3k/qoFe7TtN5
tYbHrJhVT58XVMYv8WPKOFO1f+YClrHLWObDc6dxYoOve/CFKeR1thcNQJMJNMpkzhFlDfW10H6S
nZPRyHj6TGdeGX5Z/ktmavKVmFnDZZjV4SBspGJDCCWzdyyXpgVY2x8QRFw0baFAB2toptbJo9PF
pYWSgNhpPcD2qQXxWq4eumwYembGnU1c4nTMbLMkTLRMISzPssv5w7uKO8X6IXZEZD5on/uCe2Ku
3c0fNyhr5/vo3bin0/rDPZw9i/OjNoyvv9f6ANtSM5pr/QeJA85Q9PpW/IN8VRO+OsTUvdG1eyT4
wlxCHJDk+qcHhChvM3h0Lp2tuUHFIYDXkIFbTp4xAzvbQfL945roSR+NvI/uGTQIybeMKwB/kRNi
lzDCLZwDBaZn1gjfJ1YBNXcOWpCvl0mI56iBUlCMZTRIn+Mn28SXm/m2sJ3MGlRCtIRCSMgqco2W
nQ+pMZxKr7X2wZRDe9qrCxq1GlB0ggSC4Dbhvn8tDuFvvYab53Ab66j2cgPIxKx9U3uZe5aq1JK0
AR//oxs48CezsVULW1BzUNrUWC7xHk4nRSxPnVB0rcgc0xXWmQc9aBEPFiCJ/qdfLb45ygtWXVt0
ITficz7DwL0Ay74C7EdCwxlwLHzQ0ly5j6HfsrN/e93WKHSo0evw8Rzvrb5ly84nzgTcRoPmQEAU
2lfCpvXTxFxle5NtUQb4IvRR5VKaMAkTgSxqaqLwuz9+WqUionvSNdG2pixXfScLK4qnzmWpXHXe
/Kc8Mx3w0NrXe93DerKS70Ns26MrkZkByKBKQD46eelkjGE6kYzumzt0+GmahXMG0A9Zw/TIzF6n
PrEIeC5hNxqNIAAdJpHw+f53HmH7nokd/NLaV2j71+mMpmxBGoKBsW5HbGEuZTB0JqG9FKMDN1Di
5m47ON4hfSzWMAwkgHj2keAqYWjACUfI7FfLnUkDAi4ylKb79HpqWFr02tsjuun7NCi8HTggw0+I
usSPrP9kbMWqbJI7VumQJJplYk+J0V+4tKsrMEqRuBtSXRytc75ovWJTdzv6uEwvY555+Tnqc5B4
TbCw4mFSa4uBzfob3EeeAmwjFhmDATCfWvtZG15BYV9SLVu1wmbfmI6mnT/NQBa0wwObAjP0mpTy
fC8gwY6vOfdhvpf4PXbVCwbiJ5iU8A3lc+J39NaR5qZp9GWFk3Wg0MlJcwX1NsLhmuLZixjkZtoj
QtMJPdeRLMI7pOmXl7Xpr4njnoSJ9X+w8s88YAzdeP2JCAB+oq+s3iCtTfytyqoHhxvJ52Kl/b1l
uOMuUH22RrvPvGXOkUOsEXtcXzg6zc9eB4xHu5YBQ6mOXugs3AiKgyCtXmRswm6DOaUh3+agpPcq
m8+po5qT3ZI8hPu3ATDMupIsrpZQCwssddmdm2A0t/84d9ksqUrdnq4ldJ3BMQSLiVnTQSjFiDBB
xBqTwgTOdZE7GSTyKYo3oojntydb341mCQ1qtBnYfM6zCPIbQRl+NkaxmwsqICDoE5rWYlu7kM+Y
kM/72jIKIP3d2hFPRzneiStRhMXVVRqvUftZcRhlQ4KDISvSOU6OgYfmO5FS3wJhJWjjgmUgYFKl
M5f4ASoSX7XjOMvP89V/z60USV8qS2cbeQuXoixyeU6fHTxrpClzyA2kkxJ70BhRLVZL2fk3N/dn
+WdryTfuN1e6gupxxIQ2qnszh44c+IqVP65ChO7Yj5n/7qxNrRmpxO8Wd5kDVb3ELUYEFZjHFOgl
2lmsatoDKlNnAYa7wYuxuXxbWV8AqsjEEbyw+hSn1pdB/cTaoqviqEOENOtorXItiRUP9unKZ5wT
J9tCKjoGbCECF6GbtWl3n91mLQWjTnVDbi3jMkI20HY3GCArGGfFfAFS5dmsc2H3DdwMoUd9Ygly
DFRk2/GStQ+n6QMHHRhTsj873LpO7U04gF5huzMJ+pQlGM5uKRSCed2wizlpegrS2CkJ9vFsDmQH
AO/MEt0GYR++Npe8JtrZJRc5sJU0MmGfGH57/VqjVCB+BrwjL4oKPHFFr2VEMF6WMR93n2J4ZGvx
mZrHHfos6rgPFS6/x5lMcdaAo2vMImkb9GlV2gwr0vvzHcbNSGwnMCzAlOh7NhF8d6rO0rmcygjy
EMr8OvA4ZaOLpxK27SjYrn1L9BxcmXk+/IAdnTnqGDxle+UfIcAkjnjhhLf/GgidqQPmW+++SWGw
2WpBUiBVCQdzmXalT9tdKtb2Wkj9JF7J8c4By/7v4tpLUf6kjb1PJVA66S/M1dC3FLIE/1Eo6IBD
ej2DHDft507BQCJulgZ0KsAzrYqDlHEuRwtAVC7hMiXZef3e6nA2/TZjq/XSPESt1AsxoU1Z+zUS
TsVDIJ6oP5hgFx9TdlEzOIj0h4GsL68a0NlvM3YqTyWMbgAKsOs8NMzXb/mQhOm/n9gC6f/Uj4Ih
X0ETtlCatKsyW4mbZ+YFYyZSf4utTvevY983VO/529K0jbhm+cCvrXjX3n5W23T56UcECvo/T/Hl
3z/BvMKnNgbJGljYBTbSLKZLSWvzUf4efh0Hm50OLyJ4UVGAq1+Mya6lpL3Cc46BgsE04TwsoEJC
yaC9QgHowdlxwMIMYDn4wU/HpFBMDvbtTgtvugFjyMA2Ew7fI6DVimxGQqDE5pNLpIKyjI8oO3rb
smtl0v8YAmFVwq4L8GbzuJkwk/Xl2uCjKJIAJNy+NUckkUDoonC6dpW3y9IaQZPszCLJQLw6CXU3
jWNW/wFxkWqhubDO6H8ZJ/mdjGyO3S+4bo07bPuUyFvQFvAA2yqjxie+HndLREghRRxxgaUcPQDr
AqLOUnuOlO4qVqykBl6dUsjfqnTkYxnXRq/PRFtMw3orxSpfHdmyqiDic9jC3Duo4E9mPoCretRB
9T5/qllfoBdlA4sG48N89kR8kaUpQggPZKUn36e24QOFaHau31R5GtnCTirRF93iV5slRqfKqNet
DsQx2RX1EJFG2HqquWFGGyB4z30CA+L/4NOoq2fLLvPZo94PbuwV5aw68IiCK2Wse0g6CJmIoSCV
/gvC2KaNYuTq8+HJB+YoWOVrGuZ2/3bsmuGjBKBz9mzXQAbvVS07Ei2pjd6frRzDOoltq2RvfW0r
W+t0M/CiKBBnRSEwQnhx7hfmjfkAEeZpgWgU/yi3lXkHYQ/H/culft7XaAuJ2ORWu4xY/4uwHuJV
MNZ89GCrYHIHCZyb8K/O1t+qsKCeuwyL9bDsC8M/uFMSTArGtzkEJNmHEEFEfBCIednXAzPe7tHY
YW0SlVL7uwGbgRPaJqkQri+/WEJ91y10itfndIuXs6nhyaX+8cxBEDJNMoR4+YVKVm1oiQ0kYOUp
jPCra7b5d4UtM0moSZL+9pW1ytCTz5fuP5OxdZ5i6ATnOSsSY+egJCyJjsMoNh8iFVi6vdA097Xp
YbOeqoqqH8VMRE3SRr/fkfiwJhKsfCbrIGtZNk53aaRu5aJEesLMY3OF7kJ4iGo7HY/1Y/Qwr1f5
f+GWOQTvmt/UHl3aGJAK90NacF830VWOq9LL6fBK0Bwl7tDc9Mmq24vsghqaeKciAKySbdJ+/JP2
SbDatHDKZdJTawLDnFXWQbzLLe4NQPltkyDI0UowuUTG94wDUIkh/zv33fitOGpV30hSDtRUCa6e
6F/HoPojPL8mD8BsG4SQyaSthKk6RXxYV2RlnzjrLY+WQxkCIRJaMMBwBO0s2UXhN75VuEzUvxec
8mxggXIr4NoGgfqxoIJb69XJYz9N/OnRpjHJcjMg8WCRBCbo6KNcYefxnD8nuxj/ZUFKGUrj520O
epbOBlDrD95IHJy6JFY0ADeUXJXc5nuuGZqgdQMa0hxcv9TbkrYtGMB1IC9NJaSfBb235J3t+Oui
JbmV4ZVahWJRoAxuQDknHSFNNnAhwjB9qijWSvlfnNdgAfm+a2U18egy1udWKrPr8WpQ1R+FxQJy
UiHckMtQwv8Ow6Uqv/B79aGgsuAIbOi2pSNcDz7RPNQwdWgXjcdWCtjRSR9Cy9noLwIV9o3PmIBi
vdvO8/rWI7nECGEG2qE+6uLNrRpR11R81LRm0WduZON6vJRU6SUEetcuAFPNgYjmxozRkDkHfYkb
Sb/2ETZoNj2nrQq+m2bZQdFUdwTjYdM+lFUkaaj5agtVRE7rAgqStgCNH04NuGVofMWad36WzwRC
Q1V7yQvI9aVU9U4w/nLnrdXOpKo+MjbXyc3g9+K6jKGUXuO3JZ6/1QFAVyVjlOOIPN+RIzCEEV/9
td3RTpLA/AeSDf5J+CoblFMsz/Rw2E045uPQV92Sl3ZKK+UGtEsUnR8GTZpVseElJKy0O1gt8saW
Rjs1RJsWLuQBpL/5ERTANKKCYolcn+IyGKZjCLp1l3fPMOPzJV6jsMDZXH7efwPE7yHE85sAezP3
1EnBOZigLBXoCkFK/O35KaT3/3CRTmekkPJIld5w/1zAvztuCNf6cB5ToemBddqadCCmJe4AusYV
GDcFdKTGvc4Qfl8LoqFwDVnUIRDaw/G2Dt0pnjP0/XppcBXlBOT5nCZPfaaUn0VyAhV5QFcISxy9
c3NHVpJuFdki26DWTxZsN6IXehCiKPPqDWlmIKe/Dm2DHITbRn4dLqgacMUO/65/a8+q5l+miZqp
c9yAnyJExoSFC7KinRW5NN7XJ7BUG/edKu6djXYQu7om7EtjgUGMx8mFuAqLGAEi7v3PU8rjxxfi
b7jVSFQGYcWOlSCtxtt/VmZAyvK7bp9MS66mKR0dVQLqDNA1V1mvpFaCwFOLskVu+BAVKsteTjOC
giGqxCbwXbceY1s2HZRxqKxNZfgTVgLRNpHLkOqA+fSiEToe+/Amn5USuxYbzrGP5d5oltk1lgMc
groEnwWsz9ZE4Dnxbs3eFeKPgnJGMde96a7sRnAQhymF/6inyvs2bm5PeDRavWHb7gKgK67fMWih
tdL2TRXQpv/ts9hOtCwaIqiDXUEDv9pQclpEKTcbaYq0PQnGH4EhBBgZLcepiSJ2QMJgcyHdev/m
OnAITh7jYewZ7xugJQIZbX02HwpuQSLjNcBYeHBP6eDslWEQuQDwsyzRpOqq/wsPqAWPsk/4hWBn
cOLwZ4BgHZJjn33wsCM3Wruc9dn+vbmZXtYzr+S0w31nKLMFsyyhQPGW6QVxI9nSxjcMLEEu8owA
bF25IU95BtYRpdYuRfKTmDfnt9tbesfcBmwKcf7TjmWgwN9qIZXxc6pHL9JsZ5Hpkg5OR2c3jNRf
qAXujDp/BjOKSDWXJT7EQK1nOweSxePH1yPXWm+RLrVl3Tl1dql/7aIWakuao7QJaR0MpEwyazO0
m4l1GCcBMrJlBzPDV8nyMJ4jYKkNPCuKxH6bmsybpyMp9uYm88urDzYCuXZZxeEmW7pGc9S+bGBM
B3WZcpsIwNi7jtLVB/xkPcZrYiyZ1LlEX1BfLPKWnm2Cbl8Pc51Ts+KeSVxG9wmj2BVySwcA5f3a
+lB26WO5e7gw38H//Rf+G+Y534Xv4wuBelVOoh0PrpiQ9SwyteWgwLnrS/rTdTveokMJ4mYESZSX
EDjjO2wjfSVOxkQiHY9NpCsuJkfv7RMys+m/U7aUtfB3R/KQNJ0CxH5mCAROZGNSIRzL2t3H55YJ
WdOwGNuKp/aAQNHdSt5B9BVu6TEcpsoi5W1Zm0fCpscZhvEEEvSu2/sCxnm7WVIu736Ij2uG7pSp
fR85x+jT/N9dw3Els3KnOGVnyEZpbRd5LEpFXeKDsF+B0BkOwYsExJoRROzvmd61IIlIMqM7/6Uu
1DeDKt4dO31+BNQ8S89qCRglX4cqKajuWX2IehnxaFDkaQXXGR53DrU3Jym3yEdYs6bZ7Z413+aE
0lDN+SuS8f3UXk357ZXWb5XPQ1WiK4VTMS1pu8YQ8phyVhozPBlGCGZHiQTIimNPRBmGqAG00JvH
HC4YmJ/B4pEhBeeW+F9/8n8PueND2RiX2c/GRbae9FAQ3/sCP8eg3mDg7xehFazd7RPo4BsAGZm1
mn0MJcYujrGhfLdyh09JPOOuANwaLLXEMPCayBy//IE6arxaM9K2j5AAtuJ0tMLq240A/6oSz5Uo
eqEiHd3Y0RHVv+cQ1Ueuh5ems+kZ/sJaTP3CAoefgZYewUbf0M/do/tPBpjWyFl0NeUmH/JbFeJ8
QeKWtGWLAVTpxli20Ux6IoC1KWfbl03JKUZlsxbcy3QnIJvW2s6kE5SR0ylMjfkAHenGoqclMymi
dxhBpHrb814uoYP2FpL4hzTKks8NTJRZNF06T02TRhvzpHX9mqsz6DnoEDxs7v9jC7I1pD/VWa9g
ZEmFx/8DSBv7ks4Zju2parJOWe7rB2R7+j4TvZrEB7gDzb+8JzckAjH8CgVvQrFbkRsBPirhWNVU
09EzvmC73GtBjB/vCMo9yQamWrDSvXK247Wld/n2m5HVTf1WNUev4aY9+Pffzeq8mqAAByhI1bJa
+UY4Xl/rt/lnPaqdFhXJbDByrUQLEibcHNvYET+QvQL+XxOchSNZcjooCOhz9LawDM4fe/6VFRFU
Xi+xNNZWv1AQNFtsCjiCzYa76lux/s8DcLB/x8TZClXfXrJ1PO5xj5lEwSI+4VTqiWTqG+c6Fo9B
D3H6wn3ZqVHzXU6gTW4A42kSr2ZWG+Ag+rRdysuU2VPS4cL98hAgzVXRor3LGAol/L6pJCj+sGqn
h3/SOZZp2pkc2Yjix+zv0PA/2YMH7pcha5IIUfXor/3DbOeW4QA9czr/Tb2mmjQDaea9eT0YeCuF
k1HLXPv9N/1FjgzngsrpDNy5Sy55YvV3aWBFkuoc6jdzVXJ0NULpWezahYq6rk7IzYZjgoagVpw9
yGxtTks3RY2iUS4rvjot4wlJAMdzi1yXu2phmVl3k4BRDxhftUucZQqvhsoZifWXdWCx3PrZjdFx
pjzhIRRbNX4ubTd6875BVjFiKKjaSwJFMPw8aBS8gX1Pv1m9fgRsL3VkGx3PkdQTX7+R4tu0Ahqe
KfkD6C3EuAbkb4I5wsRPgZZTyvTRBzwUxt6O4ew09cFjTE5xexQPYta0VXIKbvRDsyES/TTASw2C
W3JG+SsCZ18zKL3aZ8FwO8ZKmGdP5s5WaZ59pISYBvDgXO+8AChbTlcGp8/vDfBo7YAIb33LB1T5
KOib1TvmZE+Zvt7Ed0iQl9kcWJMNxCPUbQWZJrK8OKB+Rs+knTKIGPGORBoi4EjbFF3hf7BMCvWS
fZnwuwFygg0BKr3kmDDAFv99mZ5XJbDQt262iyJsTyboNUY1faTDX9Mt9WFXCpVD3QYDIXFGi/Kd
BSjKJyRxAfhK7g7gspgglZusABlnd3OgiVA/5T9Sd67hnzzkfmimF+QKi2ecapVNa/XoKuByawDk
DpJOagrzEediIuNG5NQZbopjCxEqG0XWV6tylREdPgNq1uaz49/zOY6QvDNt7qHSFZPMga76ItON
U6DC0gabkaGWF+1WwNu7acoqp7vmF+9PO271tSCDyk8Wv0nvM/Js0aTdwzsns4LrS+4ec6pz5gQM
n41c0lo9D8/Da5fx6Kgz7A+P3X6VdMYp1BNHpNm9f6MC5wyOBTo9eWpnRCrCgu3+DdWqpZfWqaW0
u2ynnCvHfd1Zq4D9q9s553R/cIC1Ya21OidtETM83PZ3AxQ/4lQjL4b9gqTcgOGVo9YKYVgdTzdt
3QIuHeL3Bstlx9Baai+MujGOexymVxFzFljX5PkmumfCwTltlZ1+9r+p5k36Lfb8QWMMCC8yoHiG
FMsjqsZzCPG6uC+++NUMbvc1yenfFO0Q6ZCb8xP+abuPWBIaL8AeUD3Y9c2lNUNEDe31X5OmDVUB
7SkKeWWTQDxmBn/3iyfY66aEvICdGcjAL96Dct6Ozh6VIatMyzfmNX6srEZbbfDD7XvwO/V7/4xj
aV5LHB1A/pubvrycJqsTk+ePZz1Rf7ZQaohG21ojiTHBHKoIuAu0dUGZy9VR1AjshgQ0FtKgPBp7
z1H+4AnSLtIFTH0m+Ds/dC9lwclxnIwmQPfgMLiUFZdBW2ABkI0+iFy8ZNCTI95Mww1rNjD/1zaE
NEGxo0e2t9xaylEKBvDh3GEB1pZSP2ltbdF+4+BzA10DIeUypHXd5swTbzyYvMhwE4oPAtGUPSPv
a/oHSN2xWGIH2Ml7Wl3ma0d/AXn49M1Wc4MhMX4Cj1abWp/AwhR/nI63knegPkGdOeWVoZOpZeeZ
UzqFsbTNT3TXZaSVCtl3S3Pm1nTep4iJyeQShX4agGdiGT9TV4mygltSlfJ+iaE9kF0hiTUvvj6P
OkwS1FOnqlejkAwi5PAvrrnyJrO3LX+TX3wBd8eKzAWBaBzm1Xswvac2DUxsh/unGILIbOdjy0r4
p4WAQCQbqOh9lz7qjtlTgAvN4d4x6wz2bHfoHmWMIbyMDdZdN0h71omAU3eemXGewVXMpSYGLYnF
a6j8FlghUqzrxdfoeW19cM5N/qSYY1ra7912cVYkm1AGYfnq4hLXcM/zy48uaddoateNT8zptL6A
NYqviZ9BoclFfkFJZ56UKJrynuQLPvFo8tGOUvCQQnO6PQiSLqSyPRiWPaPKhJCqah2HP5b4123V
HK/+ctwn62cj/iHgPvWd36jd2Kii2+HHNcLyu5ScJswk/PXdJ/Hjugnn8KxbjRpGEAkqmugc8bnS
W+sGEGPZA9f/g7BtvOgpX4e+9E30VHkKlPxK0VBcuFkFLogtiJ2HHqmEEpVcPM+lJbhtqYyL6FiN
8bVhE+63vv1JC9WcX0bl6MPP4sc5Lxjlk3nsh/qSpQi3DnfOq6YQwSRUugz0FmhmTEZkjMfSwGV8
hpZA+Dmv2Ul/BHp1X/YCRLv2dvWz1YDuwU0TsX4iVjZY8e/V/WWhR+KYCbzfolLmACHtR9Eh/fIq
VMjdVsiK0RwQwUIC3esv88o5fKfKHvTv0GUra5Iqep+Mg2zOvKSg17bqDQnTrSfv+QDtc5etaxcp
o6m/qTew9k8kuzkFamEZSoEjf/k0t7r5puw6PCoT3ImIUHDGRo9kg5OX0ucvb97K8Ho3I/u+Zwwa
4TQ/x4W+/O1B6ge2htVfWnrSLoOi1dt8tJ0JphNs0JbxkM/jtuAFXHoUDeAgB9Fc4gwDCxX/I0rm
n/f79IfnovYnlodqLojwGMl45qN259Bncp9uo+5vIM9xzMTTENYVWbkCspw0W0hDBVTQQOCxBGDI
yCDS9xeq1f06eSlKCQ9UzsNV833KXs5+BOruEyAp/ID7B3eSR3Rp3SX+oWkFrjxMomFkFZNNheBU
5dR1hBToVyKARwJm5g24Ddg+fS7SCyXqTiStGrxyUBz6M12EPSLPLpcxFUF32xPcVr7IWVSrYBVX
A3XZ31n6n1nGVn7Fllpsk645asWu22gTJt7qtpqrZkl0Dd8xenEK2CnPi47BL4prv4WHhbhkLaUQ
Dx+WzMdxSANDEQaVqhTUXAVDZPUXWaq8KLVH1WJQcwxbRK0it7cOwb11sKQWolWY+Rs5EHHXgNjm
tc39b6Co5vK4WhA4L+xzjxAgpmVUGgTE9+cOYfymcssq031EKG7Qt4YDgsY+Qnae9NpDf2loyhcg
GBNNc1Y5CkD5EoeQVcdI76+8QhUosoc461voFCR7liK26W69PF5art+/Yif8HpZnLGx7jo3owSRK
BVa2PXtNBX5IzWwOercRagnz7L3KC9rkfKygugQWVXiebvHUMhZflQogYvzKsDA2azg1Lsfglf+u
H/DZ1VzWmmJL3bQ64PruiTCmFHGqJr1RrtddSoFNCO9Id+CFTKJXh4IEfwk28F7xmNR1U5oZkg8H
TnUBN7+Piy2RSlc7+3TGrZ6mxSNX9Vg9jYiqJEG66YAyI7EgElv9bb8CpvOGwt9M3oPKrE+73HzV
0/rkH2sCbt9KjJc+y/wBT5y9AqWdnt2kXv/dJGl5SxNFkJNxSqjxmebU2TLRSXO+Wz+2Xc/pAqkE
o/BQzDYHSaKnPRVfK98Uqn+bHUnhY6ngCAt+qvmUfwev8NFNnCuwlj0fRfLinSvhCtaJC6A3+ZSw
xerozkMjgwDy/TAu7SIgpSKwsSQ/QI5V4mqEccZgVzBj012EDqiXxx+FCNj3Nr2bPm5e9jfW/ZbY
a4D4lOzmdUZxE++7jakWNZpV1UOhAsd+Pej8ahMPPudOlN4yFKKU4YVJosAFEMo86yrGWyeIPsgV
zj+kxmTQ6VOmeKNY8P7/5lFfa3O9q1Pdqpj6JvH5slAqK6p6uGoNVHB1Gx1fcgy2El6vc5Vw+Uw4
8tNgqhtdXRb2cOPmsok+PQf6sxFHPvF8aTHVeJetMll1Xx/jcRwAOb0qnAjKCBPRLWFdIQURJfRH
xwg2iN3RrKqbRL5rpNEG64qvXvot5uUj9r+UoPTsdMSifnhdDogsrh23rg3TSE+khqknHqgaEoLA
TnrW3dnm+KvZyg+liNM0E5FD2jOVr8HJn/nUQrKWJAvu7gai4u0lIPL1i5OgAkQ/5C/SiiCF4abi
HKQbQQ8IXUcggy4a6aDvSxwDIQvonlynBbsBpx6F4arPAUZiQ3ky9+1T+AMCmTREp7gt73HuOEBH
dGZyw1slJ20NlSmhzaK0RuOjjx7rNrf5EO5n/g3rdbZ4GzQxghE+BlPrcucI/xoX6BR7bhbajnLE
UUKpbmCnOmWk9tX2zt0wlmhb5Q62lSGpKY1GmPIxtdJwRZSW14WNOxFVAP3J6dhQdkAqUpLmtXkQ
yu0HY+Zsr3NKmTLQeEo/eXARtGWfdiFqYLAkp79ogtbdTwPFl83/dwDWXtUrhkFWf3U+cw36///o
nV2h+2ZAcvT+H2lTy7YiISF+14MR/qB8rY4N74/tCIh530kfheariLNe3k3+aOZ/yrIO3A1tjojV
VqTwaiOHCoYRPeNZXi3GQvQfGiJX705sU8YZiCVsnWBXV1lXqe7nmsuE3EU4yfx1OfHPOQiWgjGo
OXoKtzOzg/3WrvEWpA8LI0z7xj24k7hxR/aLXCz+bJYM+CnsYrLi2TaIz8S/Xx+VlAbrnU2xxTu1
wok5WgiIToLzvHFOercJg8LjNNxRh2cOTLf8iFbVY6GTsrJBXHL6BemORsaSCnZLS9O5r9LIjJFV
Wa+2Y6Zpa0NhamLErKVIqlRjZTriTVYqZsdQWLkS8h2OnoYgz4A+uNoWFqX9Q9CVwFseiklyk7yj
dhYOXGXCk8dmDFRC6pZXFUVAS9Ac3kn0C5GodTykecH+sucRw3wje0OuIyNWkphNyxuAbPLZnvCA
0pwQc1Nle7HvLbUdokhNeNEJ1pKXCyqZmpSni12got7QcGfyp/euBnVozjD2zLueK8Gf7+Imkqxm
Ypj4QRV9WQgzcvgKxEIoYwVr9PdyMOxTIUBQ4UzTgV4LJ+CWXYh7djVT7CnDxp6K3ZOvljg9e1AI
NeRehMgL3xop7OD3yKHibqgylANJZ/BvpCaVYBk6qkN8HlWVE6QTGGUrZV0Ju7B83R5/IuEaFkiu
u5l2wI8bYtNE+7ZIiO+0Q4terKhwHSmx9HYQhuHsqRrOFydQXuu6wE9TO0yXk+kO051UuCbQAvRH
FFcZqYiOujea8EQGbPG/gqe0yygj/iarSsvJgagiE0qX6qvhEod/Ximd3BcyNYXH2qkczAE8LXwx
ki7uCaN9U/DK9Qy1iLl3aYOhYaYc3ExpjjAvFQF9PIr1EnVq9PYs4qxqNfUPjajy8BjFR4K1fSWa
e9ouUi4+T/eSiePQOboqTUThT/KOvSh7gAvEkJ6PcQA7CBwk15MhfhJ6K/M5s1yZguJXGLhhJPBd
VZszvVRHcBM//upurjjuWkN969hxc4xLS/K7Z4q5w0p0oM1tt8NdDyac7lEa3m6waw2aWjSbP+Z2
C8tObsVLtWS0W4/jmZlMlejNrs3SR1cxPcZMEYNazzQN0XOOakER/ISD9Ekx9IgNWgVdtEWxrdDh
B1GIXlLOuJWFEWjCuyB1IL73ZFp87yGiLbHdyDg/4BLtRfm1UZMF3dW+1fwFDc2WmO96W+QnTVLt
N9WHXE9YJdwEWLj1WDU/5eM7ZzQhbRaKFrgFaGF8kyEI6jE7O5tAjD2DhITTkidSOCDFPyaP7WlY
O3q68SWy0sR82HJ7ScriWe/vQcT9IqJoRcupFDwkzgIoGlF4DecZ5qb5Qy2Jxanoba1QhyVjvK2l
755BpMPYarQh5GCbsRzzzpIh8wfRa7agAHVwpPXi7MPK4hy+CT17ze8a9fyKmwSuk5I54EgZSgCq
FWY86MpKlMW9kB0A/JrLvZleR4yqfAgnMnhRJOejVvzQZ4rkXujkc4Yz/mBUGF6+lnuWqXr8GnBb
4nUpyqL1cwPSMBEY+WUa3j0dvlYJR24wb10mAL5vNX2J3QTJMFcmBHvXL/5F0yHfzd7iLmfgzlkj
CVkBWLPTQej4l1Ud3aKzi7ib4xAAyPr+F35stjHmG70F2zoSgevnswb7U2pykvnvVYvnz9RyZ+9g
56x4PhbPd5zzd+uPZqqZrQnKQ1e9kV8dSZq40CGG8Mlh2rhP0oTHwO/uNqfJ/Ggvfs9+1Y6NON29
wr/utkI2B59WkZcodc4cSAPSpWYQXeakLmBgMZVst5Zlp1OgHeoRvj7xnHh8Dp5e56Rt0Tss/+5D
qyehAgUPX+qIEJyBNe8AcHHccDBgcN1zGXCQJzLhe3DlV2EVtmtgB7Lz2IiFlslb3522pI+busjh
YRBtHt1X18Yle5cn0Zp4KQ899Kk+3uYyFp74K71EBMXkOsCR8XhfMm0FJr1KgJlyvDZheT7W8SJx
Wov2H1ab9QuLsVKOdWD9cnJNF7mgjYoe8OMRy6j75o/k8MkcFykL65fhzKM8TxkN380qyW3bP78K
H/i6nFC6JUpD/yMUtIAOFXottInHCdPUUAmbEuX/GtnemFovoCE99Hqc8n91yD3vjg66ZFa9oTQP
xVb71I8c+QtUwi1f6DzWvi4i50UvH0cLXd/iLY66lRe1x0k9RRaEdCiklZb3DZkSHmaxmNJmmo0p
b2haAKE0KWwl1W3rTkwrYYXcmzHqwRtkyeIB68/UFk1niiEF5pDC1r3zDNg0OqimiF2trHNqQ6Es
i0Mm/QB56NaKWhhIPPi4kU9eFB/ksk9PnZSR5wsvukwFPlfHKBytvnP6nAv7eaSguyMgiHz2GLZE
vPMHYpu7yFizKmX/89avXfuKEwuaOR0r4bcUQXY/Bc9mB9ZABcceWquVv/nlbXtM1Q0hyTe6deXJ
r0AMEpYefyvSI0E4Y2j5I/gHDEhWKJC/GCQGPr++wtGMcDRWUpqd03OlJ8gorSoXOkLHOqN8AVHW
uRQcV+wJYPlBV3YnelXUgFO+UGwn39yM+ATuwC9DnX65YaI5tk6tG6C4ZizUqmBaHKRkrOQHX/76
HiO9WWHhEj+PUO5vbKZdfqtrhQyOVSJaH2XV9341+4L8TG6L81rVW9bUZZEt0R/OrbGx5etprHLt
VL8BCX2u5w0/YpTXkSoNS8xRw6mBAzPtT0/szbJNIqcQGMa72ZOeWkSsLgnTutpOXIMP0Rwysel/
ApqW886HE2lwK1Ro0sLonr4Dw1n4QsND1hA2Grv3LODmUuWlwdPuZVS/YlAVvYV7sga0/g6wRFR8
K2g4ScS9fuOnYztTaOTRPOTVW1wUOQbg2yxFAQSte6qbBs9/iv+AS0aLU/1gcKwsfRmr7MD5Idsd
tPlRzKRf4LGX0wC6YUOKN9GpTzh6K62aWEA6IEpcus42B9Cd7DtXSwirj09kDLVc8z/DE5+5hGos
hpyZdQ/CqyrWxLJbzCojaBtmtgtZRS21jM7qFYFmY0B49YHAmbwf0kzfOAVU78qZZyLVrkWIeEtz
pxNFpedEYkZEVD6zFla5Sxkvk4u9N0/bucTAsPmAGbhtvfQW+DxsPsF3S8/hODu7RDb0OU7b48Ra
1yIRRNcH8S3MQjFo6f7FU0KWkMypEYi4htPCebBr6S4oxtEqFDwOR+ScgEnBwTfkQ6GLN9T/b3r9
+s++fV3ZpIeKgUX9rIWjXRrzIGlNysB0LQgzmRbNjkuWtbxwUaV7594cm/D5boC9k1hYUesgCbUx
vXh7DxKcJ+a4bSjYAsNORxLHL2v8rvXlMG2BHsWBe0W8SJJXBrdPcgEAug78rRYzVZV65Mi1hjQY
JFLa73TaxVk12aeV0+OeXpuKKPDy7o1feXJDLEEqQ53lnUXdRXN8S/JgGcMCXTmK0lkxkBg14uRl
M78XvIslNmHANy/+x99EYgCa23VQ6FZrxDiZ+sLLvNAj9fjAag0WKMwuYq8WAkMGAWosCABAPwzT
sDmQWiqNlYmEv9ZONoL2xxJRfD1zGK3QtsXABViFVuD4VGwgI0ALAZ3aihjAQcfk5wxYFdOwmK8n
K5pPAnhgGOOKBGbXOLKQkmo68pI5+9Bb08JM52KOf30+qRYqjT8mwOEeuzvBH3KvgOeOckdsaXdG
oatXuz+yGXXSNtJvTPe6DtD9i7iVkLJiNUH1zFpC44WjL51vn5ydZnJcntDWa4j9MHA2gdAywOTh
ACCoIS9hkLDD/5ly0ptOyREHPbHZz1iy5J8pjddcwPjNbnDGKchQuE0J9xmei59UjZJP+vnHTomQ
Cw4Wy+Xi3H2JO92RCjMvH5ejtYUwE7z6X8ux9nD/XSW9myqwN5worL3v1nXxDzU9gDanPObYxruG
8WAeY/g7SwRMqTrrRyK+sXywgZyJeqgRIRGKpAEEMihTmluau91jjpKSZJXLBVRUQSNtpCspG/Jr
8piPmBIe7OipVAV0V9GoLTt2RkOXUuiNFWalbE4ibocQQ8Kwm5wXdMOpA8BFmGMww3ri0WEo3aSh
yvr6jnSIB/KR4YudUf6Svs8oHJx4aMtDbGzt6Kv2SlqAt+LejyUORiY5tX9eRWLZ2jrsyZ/WfmZz
iiq6k+i5CjZwDLoiZrTOncVReekF7+NYNsnqSvllmxHemQ+/vJSNxPxPw99aqODpTpo8Y8XegCsl
+lIIY3ZWVGJdVjrrRxmWPfF98MOyv8chCbmT+1HZZlXmFAAqIELZd1I4W/NVOhX0wC3c3O1lpnAC
enGgOfWoDY9B+3RHYXSTvlRkioOa1ztOOvtBF534AnB6j3mshZIC4FwVewS2oexs6trEX4bedjsC
6jjyW4RAvi63HXsGHL3Y16EjeGY5u6c5XQ4mSnEtUmsKAxLgKj7rPWMAPsKIMYVOncicEDaLChYI
pKBFrZ2ppCN2gbRJD/K5Fw3qkTqOKVpuwWhQ3ENpbaftgp7Lv1HZXr8nLUUfujcKV/LIz4ObqX1P
jmN5wrDydpCAHXpfVfcRUPGr6je0CUMJjeK3KtOFmD0iN2klCiU/JlYcfFmml/b5fCM7IhUrZTCT
kPCnqB2pf5KNgpmDxuyXovIfvCFqEF6lzXen8TRfuGbO649Eq+FHKXeEJ61lisyCi/ju36xDz4Nc
Zq4CzTRXfU0V1fQJRGJ3FpZbHcURkox/8m1/Nc18mDw0teFu4gz0avloGmJd6dn2qyyE6XxjV5TX
qzB9nXs7/Kds/e0a6itGIlh4zUUqAMBU4yW57ESYvspc1oSa3dhEgmHiRmVYWJHy+8SgqP9dvTwp
OH7vEIzT4hHaSjJdB3LTqDnWulq2/f3ME3WhxkgZLowVzLqn7iTcaLXbMw/7mVxFoXcgszFuRqY4
DlhlsFINi+EmLVeUC+brLQVuoF76hotR7jbaVarl853jduCChiOb6H906Iv8kQRko0p2xYCrgj38
XbdHbNVWKoPgZw29qN6FUmNTS8jFt0UaG80pEemxvryynH7AYLZJmGmT0tH+RJMvRKu4qfGLKoyf
N8MD9bW8j3pZYXvGPgraCP6QuDO0kr81rbUVqoA+LjSRAaxWIAsMCDZvB+JlsZM96YgqwiOHE4ZY
FKaMbEYBJKHoSjKvjzqGFkyJDFL2ouoPNaAHaC+ukCsVScWfWTHuOsQrWFAeTTgpVwhkhnMGy3Tb
sarHEzI7J/bYEFO2WEP8XGAtEeboUlf2lDoLcV+6SHUCpTMpjc9A11YR1+dkBbMq99Dzx4pzxhgP
gVPIblCJPufjEkkpZDuM1QTf77EOb8tcdQ8lGDpLoi576nf9XcBlsQO15IVpNk3VRhTRO1PUhrxa
JoSIZ3qPkU2rIN51+H4tm5b7R3JbxL7lJ2KnOxianlyE6s63xNDIx0wKbJ8I9FiS8+0i1PoP8kDW
SS+HaDRG+1zn+v5crVpPITsdbcVugVogO6qHL3SghD6Va2VeM00G0rfgOolsAySulXH1zuYzMpCj
JnpgqQzniUlYkk1so9PyXikGaNZMV1fPS4XzKx5yTbAaqGjG0Y5EbQvaVp0SHI1WMHo81ICiL774
TLl54G8gwivn46YIvIxyc0d/5pV0vFTmlKmD2kCpYCT0ybjKdLrOPS/2sj8oBfzl3ZELeMygt89U
QXqiLMp5Cngwd7HsU6/uR2YBFqnWMhCU2evL3vgClocFvpFDuN192RbcXqUoQMohSU/b6GuhGFmW
zlSK4n1r9cO/m5ksZHksXOXgMAYu9uGv3WG7qfLerqWoaByAJogB4zmvoOfOWYXW8cjVi2RcZz69
2UaO0RWXGJt6IW2d8cvyKOwaYzy8P85rvTpsNoV5x6PrCasY6uDSxnhoLr6WmZrcaT1bSsZPfBG/
nQgTJU0tGd3hEtujOJxMZLwEoU1x99SSb4SvVr1retdtOggNWvTMR6bDk0H2d4EsyKniHpN5XCv2
j89lE8b93XJDUiWYlPSPjn78UEh86X290gP1yZIem1BGm7ynm2woh5aSvL3aueKfdiE/Mmp1w0ev
uK8GBZDUGaHfTOwAhBoVtDbEgD/cwgzWecSHVDOjO+76BOWbjuJ+uviY/TqKeHr8SbseIQlvZqRn
RsAhh4lAIMUFZD4iUD/12IyA5VSjx8vyxA3lEP2PvHLBSjuQRTdW2LXUP89O+uUfSnO4Dqk33Ctr
ZG+pMbY24FTt41UT8GHnihTIOdSRjp1/VgNn9g1x/jB2RTTkb4mr5WwIiHunFLQMnP4CCkXCRGWm
MbqvaFaVkXkiXQ3pzmvbrrBJ+zPLo7hdRRsecYZLrnJv+W8/IdRknih1/DdZ+gd5z6JXNhU75SFQ
Z4wLZJ3ESbqPtzcMKZ0Wp1UXTAoF1bi3qDGblsdiy4XaiPfaNS5LNy3/7r5Rbnwc9P9M5Qf4JTTD
I0RWPGSS4jKUDNVvsBY90T+f8v1lPKZizB6JTzHt7b+VJ7/YjioZ1QsHct1Wi8ZVAfTKJObvqKu2
Wqy0S20ID4tF2sLj6L0Q+4w3NmXX4Zp/fqOE/81k+w0BuPLqB1z0mDdtzKBAVbOrPuCE11Wu3fNO
OQYvD2Mdu1Qq94lQXeXY5oXMS50WzepK1Ef11FxQ/o7fA0IJdlmUwQHGncCTBvt+RpKXACaop17L
U9v740cevoTWF4L52e/2OJtKlCTmxA8IEJ0Yx7MvGw/Tb9Hxp4j8sDt6oRZf+ihlrzVGZhnPbsWR
3HN7EX6o/x7IaN6HWnDyH+uoM9/m4odR8npPHZMTOHBNaw2dHaQnrqUoJF/YVEJv5qAiLeeKZAWw
4owY8Dq7jh1OrNDv0oz56dpox07kdn2rwq5cXvt4PWVhM55p/+r7Y7g50xB4e60nTYt5MWQxPaSw
6Lf8dtpO3mgYlRg0wq3Bbgj4VNha81seE81QAj1A5QvhdGjdUVQb1DdVSqjIkGmFwnYB1xSmTNxg
yYOtTmgvFbTD+7nSFv045fJSN8cLluzgfmN4IuwlaqAy9bo7g760MvsvWW2F1ZdzGpe26NzVSOOC
46yScttel2o2XUmZxRLHQMoYbV1GeKP7G5Q574FjMfAGmI0sX4VkgSW9lA6btVnKMvVNOX9QuqMd
LWk+uCAdPzmY1ac8sAUgFzOh2MKGdTKaNSxUjJul09nM236yNaHpqLdoWOx+2tIbLtXIB4SCie+k
kcW4SnaL25ySs01lFF39LfOZAtLMZCP/DFmZ3Xebec0XvCQgT0QFI+X0rxA2XjsCEe0xB0o3fpSK
NofYTwu7rNBzGBSbsEmsf9zYuddWT5e7jJeE2WLS0HljuA07pe0HFXZPGZl7YXTZ2lDYPW8SvjBb
cDNGVaW8Na9YGDJhPfn+r4nQQ6Rly3Hrk1GYUVJ89bKRt/+cBC/E0q1k2OXhnqcduLEAoTtBxT5W
Z4XZORCc9bJJtFPFumQfq7dXHCE+EZxURD7+hQ3Pqb+8ibFg3/A/7GAKEVo4Pn5QTbA00keUdWj9
nRdKHN7Y0ikF6N/8YQs/wboX+HdLzdYl7nw+uPLEz8sai2tUZpFwUECmrIbiDMV1MwY/m4aoN41g
XA1eGsl2tEkfNURjgDsi48isbGaUPswbvTwBbAxq/KWi+UjyK6UYbwd/UB4WgyyA9zH+L9KCzbud
mqqtLrdI/B2ShpwgJTbAdmfH0rxfp49GOcIwBOXzNyMl8ydFqMj97jvuh1h1d81Yg5CphuPixew5
vw9tRNTScfjo4Am/YTp/SqmUIV1dYUPfx6oTDOWNpbBCJdiL3RPn14+nkRGuafe41ESqIHIk2/wQ
uAERaBMbUL0iR5ShTTOLsx84VwiJj55O0stm2izDLm8rw+t/yoIx4RUXzY36+tDdC+F3IZfVu2n6
PwLu8usRPbRA0gAVAYzIVyvQkMvwBpH7ulg19arp8JE4Bos21KwTo+jnBxBJj8L7x+lS6j9Qw9n8
jypa7P0geEkQsNcE1Ny3+M+K/kImKEplgj9Ss2OAIN/C6cqLFf/KPDCjrkuVlxkMPA3JeG3puhFu
BpkkIR96w+sYGkHnY72bKQhX31SL4HM3EcPnunL9GfhNvzXk4Sl3aLVtxaI8Pq2rq9E3Aa/+ice7
29FI44fjzpSzs50Gt/2kdV1tuG+hgPMTWu8KrQdXIuDz9KtLEpsdXmREwixXulwMv5R//Igw8sYN
DBbUfuGGeUVS3jjTxdm5e5Z2cWb6RXEXU5QVnGyEpFOrKb99eeQcs82KVwNZcRntpL7/hPCl4/0s
O/bm/AatH76Mmn/kDEuDBukeVpljb+EGarSg2TbTfR5SeIfzqY0HmTjYJAw+uHQHSpotzUgyQUDw
358pKKeGmIv6r3slImraOG/osSPRwdclOx5aYPV3cwDi1QeAoD3egWvmo1tej58qL2BxH6CDbc/V
Iog2C1ysTJwDZO54gfJuGzThdtH3bFbaS8DPyJY1xdVkeaURdc3eT9hicF2ZzjXn6bOVzjikptkm
lTiTKVIMjb+ML9MImNzLdPDvwx6tKKDZJYaOu3KuIpArbOo6d5F2QbGyqr29yVUY++zGMN6OOiUc
7ozPdEC68KKWMNXm7vzunQI1AVPsjWRh//TNCc9oaS03ojCUdeLjtHaAqB6mSoVTQEjtFgjIM4MW
3bDzPL4RCwHrIXeQILlY4WiGXrS12T1X3P7VzZj+uk1cpeFY+snm9mm02sCerMkC4B/hHa4MzkjC
j9FCjdSmuZ6sBu2cNSgXBl56szZOQ4LnyK851Rg+9Mj67Y0FGvkHsomnQaLQZCeIcVVG388HC25/
4kPlS5s5Yj6vcoWj8Jt3MpQgtrsL1LOmd4VcoZudk7leqrLlAjAXei/gc8ZeCTnJAsnnbD+J+pO4
SmdvpF/fznT6uWT8MslPCMdhre/qVxIAvrum2YUMCqcnCst7TwH8RWm9+YR1AoDvGwamyCnwSyrE
DOTq1iUuIAjmU5qypP7SSXp9KoIqS8+NxfA7ozg7ihSLlvLkppAzUnk/0/Nomb63pBdRkfe7YA4Y
6jQvyfYb9mUK2FjGhCQD2DVgpaDtnqMh1PYgkOjhJ+qd7C2pDswBCQx6E+WyhQLs0M9eePBiHLoL
Zy57hkEGeWYi+qfNfXjnl9vhHjSQjEctrsUCvFQWIPqzb1Fwg7yJHYkl1IrydzC7BG1Ny4DdSoI9
vUrHvaY5CgObYJ2thPzregqwl38hY0pz6fiSL6r9OIKpSm0sLcTBO64qoa445vKy7EQNC8edQo2F
M8RC2kMYY3ZffGVfdV82vT3AJVHYs6It2d13lvQbuCmQS7pkgSxEbPc2JfYAKyb80W4VwChTnqbv
OEXQ4ysr6buTLBj0yl6DUE0r8YoIF5r8FBWQPNIDkEQXNF0eVB79/b+u6t+PMIv65T9nGaGQnEJG
KHp43OTbZHx32DL0oH1wN/YcEg9dFCg+dQqQ1QSNKFyxrmeKxbnv+nPvdGy1AXbVbQWcPAXUFI2m
2qH8UjbVI/Uu5Ls8eHk4fJRLop4xC863MaF5tpHdB0shYUuZvtRVG3gKr1nqYeHL1kW4LLmZ+uVh
V+LNz9J2S2otQPBxzeANtFeZ4mjS9nMWW/mZdPb7Y7ZmiRrjeV6z+QUrECUBO5kzBPefRMhq8QY4
p3nsudwHTQkbn0R9OY4pUcrqnlPFiQ3FrOjVb4vmekURelVtFKBdM6pJS1ifFhtj6PO8jl0qnaeN
EZy2njkJpmwiYZrdOATOzZEnxNxrWg6CvEHgVyu50YjUKwT6o3jg5bcDzP/N6qA4jeZH+fZgBUJY
RA5e9hp2BpJ0k5U+/aClQr/fgyoF3llCw3yr6+fx9YL0XcbN7fGaWnnfJDxU+lPx84b+3iXXscIZ
4tZHizKj9n3L7c8ZPgx4NfUqndOY7C9Qb0a4igj5qx7ujY2gOllgtRFbivy+39vUy/6XAngPkJUi
CYg8HwGqxLWW8uJLRDG9R+zCFRF6ohZySDsohnNwMkp7mxKCrGexwi9V2R1Nl1cJjC1DjjcMlriZ
XAw9Sqoecd39dq4VAFm/vecB+dDS06aQ5mYW4kphw0BsyYC3lOKfygn8qnxdK8h3YlnJUa78S6Ll
MxDRf1voJ1y4ziNjDiF1+rKMTK2IaAWvN2kwqblZaVUb89vs6Opn8GXEJH72APq0hbkA63ogDOeX
hnCXroDRkxH0lHLQ4EiHWJEzAZQruJBayvm+hWiIC9CAfPJg5FPiQvCTZCvGUd3qU6sxMKCqeKL7
PmQkrRXmw8Z7vJdLiRehZ2ClFQf1/wI14PPKNE8O7o6N/G5Pto/ZvDM5ofi9vscQw4yLbmOycREK
sEp2E0eywgFHXDhFOHbpPP1/sR+GdCPxD3GN8K8O6VSloVpnttmOUcFp/vNkXJUhBO86q+4e5F/U
p8fgk5b0mDb4TUksCxOMaz3XnsVcJ7gPMWBkArXKvyABEKo0WkyhJMsd3ohvwG85ZIufYEdmx+81
noWh9WV8eWww8x03Gj23dI7TyrBZxiIUSeQVycSkik2Ywk3E3SpvkbsjgyHTRNSVAuzKIHIBZehh
jp7NQdVbIPKpya+GIIaHj7va+q9s2P5PAMHlJWgJwAsgZshYvxBTniAIc1CgLR5jDPDInsTVzON/
rcTReTPN+xhf4g+xwZSE2nYByExlbR/+UJJV/GiJ+fOIEB7l9Ir99JZGz5js/iKVe/vwYq70Fp/6
q7A6e4ZM9ijF8MoVL4Gvm4CX9SrHmRjaDfz4F3mMqznGZQiaepYc0m1gTDOmEV3NKTtd2rFkhJsg
zfe31X3xCcfbupK5sucJZeYxdCBw4UaEsn+wlTIUnKC9WTIJPhjxWoKFhMiKasbxY8eE8zk0Bgqh
jMBBXmdopfk+vy4vU0D9xAyrjUPEH4cy7QfJhyhqGg75PEnS4DzS7KX4zs9jrNDXTPmB8t3Ij2hc
VRLpnDhPNHJFQ/JSNf1AjlGuUQjD9pxnbK+z9AAT/bZa20WXzOFLg5BY9fEKeEFTWXe8kSYt1zBV
1DRGtoDQN2o/ucV/imbX8k9EgQG4Ht83e1Lu5jHnvTYa7bnREIIsenEgZdOB4lALC4US209lJNK5
3dr2xrvlMAN4/Dqi9A/vJf3shGhAZ2btvMODRFQID5cysTeWcNNgGp4f3+LJTHu3GxlshQvjYpvc
qhautX9goUIUFqyXj3qZykXxtB0xbYyQc1HnpHtC68bITWIIdwAzEEFGQcs2UvB091E9Eo0TFiHO
5kxZfDgf11KuHxh/VfkJ379LkVa9o8QaAtmfchwGK1+HLReq4QcwxkHMVNga9F6BNQC/LsautGu9
6E9OFEknkQLIs/DdSsX6YXkI5GVWiFH++lX/5htheGeuho49z1NWd+SNgoJ0+9x+dHe2uc+Uy+SD
a5UUe6OhMLiYkGkSgtr+0NlnUnkzhAx05QRzISGF+SVAHxrjUQtnkvoZktrOEQCTaGS1aTVWIqNN
6iM3gHydQr7y/0EIp9lTJS6menrQpfuV+s0BGaqW0e0OWXLrcjNlAFhZI04Y+AUBMbvgvyuvD8qw
7fMKLQo0Ow7GkEw1fOHqoojtv7pgVRFC3VNH2nYU9Pb1CtKhURCT3bksBvGAthPP+VCAqURZLt4k
5VsIHk4gJ3GXMh9X4Q4Oy6Q88qXxGrg5R2LhB+xhdv/pqNK2WWmPci47asPWXkGPruqo7SqfqRWh
L1DODh4H60rwxlooCT73WdPt1f23eZ6eJOKZeImszQCabmCef7zkjao64vAKzb7rA1n9LrtEqvXS
u2gi4MKvPk8piYQlmNTFiwm2Dier5xXkntxHtVOTHKnQXuEYbilkbju0wZk1xdPJExsNfoDwYkB/
qxJvrGAUof+Uoi8mTTciAkSSFfTgUI5rbnTlbky0pStDKkjkXeQGAII0hp+GizTT98ndxqI2KDck
ym0t7UBYFPJJEqNf9W7oAP9VK0lxIdKjt3Nm0S/9WHt8iPCf2SpbXYUmq2He21vqJubXh1usU8O3
HXM7lm97exEMcsbhCSBepG3g53zThn4ZmfS8/D197C6RPuYf3Thi5K/VQkMJlXM31FBhTfxt7yDY
Vrkr6QvowMvfwrmiV+ru+mkNgvyq2cBfLnnCM79t3H+yo8C5/hnjfC+nBTMKQXAoqfZ+sbp887T7
X8jh6h2fNTmAbPyEKT4QoirY2aqIGoLp+VM99mGodd8mc52IEFcE6TGzlIFqipjZ8RTomt7gSu18
B18H+tyn004H7LsJEictS5Jj/0iNg1t6oYC6emO9XAIX/tpYVrOytH1VI3cnXiWWc+PIaD8r4tXU
5Zn5vGTgKEgG36zTzcrUflE9ve1PByJTwqr66WuSsSlupsF94+560QA8lRtZVjuGKi3GPBBNFgHU
ABVXQVSUmbFlSIHTdbdhCqHZg4OCnMulBUcS4gDlt07Uzc68wFcUhKNLzlfUZisN3Qyaxc63DUdO
oT7JNI3sFTOGRAwHr6C5el8oKL7i0tC9jhFtvXrJoGRP/gy8qsPPGRcLmjzmY0g8l8S8O8DmCtBB
YescMNHy8tZ0/3eM0Q1HWpvQr3Cc+4juMnhnb8KsJEOu8/B+mGh627TSDVgTqDsHRi9/Fw+GRa83
XWc8eLKq+HaeDmEYi83WU0EDb1neqE1QDHQs5Jcxp8Fsl9TA+tTvFpqczHY9gmGHNIZ7hMlawLaq
+FrM1JPbqPdN7Wr0e57fm8hDjjcMEXeNa8cRnzcrkGUwF6Ofn2TyMY5Pl4QTYmZSfm4j0z3Y0ZVn
R9dYWvnuVSr7sza78awlLOoiwSCwGWzi4f2piI9BVvDh9YFjIrua0lkfX5GYUal9JAmnO7i/U2qX
klFldNQfasBthYSxeou7uO1lhILmWNcgwBERlwhm8Q5zJGZKyAja37eohLyK5of6f6O42kto2MB4
FpDyDVWfMoPf4NoZ3qB8F2HTVKFtougieqCWeKuKfaBQghTwAi7ePBqyd/TF3zjayH6L90h9zfAG
iODRCOtHq61SABTjPiPyWE0LpwpH37L3a0A5xYIGBdvp9kPiVW8Db33+QGGncXGXS+bad7c/PKh/
fQWelQtt3auB+z794mlsEZ45anc2ZxcJpcS+oTsHEg9f8jn2othG1CeUSkx2QL410BvP0iTExekv
cwUBElUUmvZwo9P+/XXy6c3uR629uDJFN8+uhDJ00VjAAWjgB6t2x2OgRfnYd6SURre//L3Py5mG
4piXsuzNDvRCDgf659FbgcYCcD6k2yrcD04jIF0Ymec6E8D77V5d9KuXM9n0A40VVa47+WBuxTLc
KO0nMZBNUOU4pxhYodyVFN+RyGkbFlZQKhxJbXsvADKmN15NZK6md2UIS9wtQKS0tUepb1xhN4mY
ucPzknE1ycsIgGJayIIiNTAQn0jZaBuqsVtph0iNm2rpnQc/AZKIKLQEJAR0lzPqWb77BCFg1yam
pco8icN1nRSqVghtjuA7X9ooRtloOTovBMMib03OJ3jSTHeorzYEMizX5tPXKv6cWObxZY191jKD
lmzic4SvM2HXGtjqt4UBy5dHuYtg5VSj1+XRMqzABFrFj+KxqC+se5lNgTyeiShvBEY/iMYhC7fi
2gga0h4xFLTTBNMlKhCwkZsj/KQUbBWMmtbv8Uwzfgt10imWs2hdbmtQz3mWfHgO9b9tUdYMvXrW
A+5y7WranNl3gS787bVe9vL7PIkAF9q5m0E8xb/+vtEMsxdXedxyuq7zzJwjuwSo4cG3wNjF14pf
aCf+b+oFIWQs68Qit1+5s+K3M96dyUJuKTXwgji5kQCTy9iRkzOEBudV/+Yoo0mf1Khewp8MeevB
Io5FkwNk1+Wp9adc97b/csSvustu0QJDHtX2p4ztqXuFPc004tuCjEOSPUipSD75trkkq6F0Xt6d
o5ZvTU1WDo3cmJ3oZMNN+doGxcVo5/35rB2/XZTXuugjfjGjlL5UwmK4tcd4TxWTJwMy06aq4S1Y
vlO3Q+u8GvS5bizRBqTgnnnsUkF+9mldTAH0TVmSVB5ocyb10FqDLZXhwdzrhQbDPbQ7nlDto5Kj
ghAIAozBauJ6gh2N3mXMFTEQY0cMRdjvI381nPfL5AdBAHVw4XFJDOy/eMN0+oaZWVIC0zKXHDQ/
7kkJzG8fa1lcK2s8cJaSUgIgWySZwuZeVy0sV24kafvGQiOGVGpvusKsQAlDMMeSpPiHFAqveucO
f7Sbd2kP9XUj69PCVbgd7r9TXWT7fsyDz2BdQf2W/2qu24PXB//DRtQ0U0Kcl95yJEd9A7HYrHUX
ZuS1tjpA5tw7e7Hj/FkOj6yI1DwYryepSIT7B9c9X9WYrVskSRRlCQPL0TugJWTwEKSyn8vH/WUP
AlHG3NoXjGOXXAy9x5MGthWr+5QCE8n6lh1g0bmytacPELn2EkaIHVmTA/AeewF7mwTAfINIU7Wv
G2qs302+eqUdOtqOt6DSxbUL7WdqnXnUd8fio1wgKuvE+sQFidQynIVslITJV9XW/WpPss1UEmcX
MyGnhokV4lN5a77+UxS0+n6/lHe/ZRMs12aqRenHiwvyIH3ydDkjQ+qGXu2iYVnFOg9Y5ASBbvzl
m0nwAlQJ5euvnk2KwQ5sGnfCpdU7e9lIZo0VAzx+n1tYbM+olUsbYDHdiTgQmKYQH68zH5afjsJI
DweRxhRDQJt2Pg6DgPYpWJrrT3oD2jJLy39ZOgYeZULSwdg51zsBBEOYMkr4o+0sOC8HFJXOKEus
vbDrNxoL6EGL5JPrwmez3jqvZWreSKNSDiB/svSeGMvubP1gtUEd47DLpXedIeAL7Pv5V1dVYXHg
b5+RnPT3RmyS70kgsfW+H8hAcsXipqs2E8WCv/qJGk4Om0LKtmk8p5/cLeNrD8PJBb3/32ghuIDJ
Y9Y0j+9kMLQ+sLKjSXYjeWBvX7NB7gZ7jxab3pxItDlK3j8SjAN1im6Enz+lRs+0GB8ur9ispNQG
kzJjQwOyB5SWlGnz2sVLzjwOUbC8BQuuR96avPo7fsh9TD9JPvz2sGgBniHUOONHA8RvGNSN7Bo8
00du241Z2jREaNaKxsC7lnvOQG0idE+x8KOZYq/L7HZe+JSiGef7C151JPYAWabyaYtvgRtTd/iu
epMTBsZkDc/ps7DKR5h8LZmwnsRJ7UEBnthPC4KlUGmoXdayz+kRIU+pyXBhG6r4wbJq+yCqn2oV
VUIsuLO2uVtHmboEPNcIFJq8NrZrie+KqgApipfqkqMun2fmN0nvhmkhIFFIx2jMaMkAWxuMBCIH
0a45C19G2rlF2oIkZndnAr/KtyxlSIiteOxQOv++7ikanYwVrhkfBR8DzzFCb6ejePvEs5zYad5w
Xy4kpr5fcRo/wbz7lXFVaZYzTd+zweCniETB5qsnYopfqGuoN+nIRT+p7DUvC44Lg9d88t032CL5
oZj7NmDWTDshOdrw5Us0fB25fl2lN5ArxPqvHsN6TMmFsqhh7rvLax5P2tEp8ciOf11le7jOSlhl
0Nma70A4CR0D5ZvoFt9qy1S+yBl551ZniRG3pR/DfD7ND/4ZpG+twMUFNkACkx5EjW3Bdy51lj4e
wa8VpXY1ZWMYsZAvRf34HV/XdaYVQYofA4W9pkV1VWK2eXXauQAAFPEsY1PltF0F0JeYzmPGU6Hc
6fL+TbYP4ZbgWYP9N3Yxs/W6B5FGVIJ4rpGVnz7f/LbXTWcoqisRylrpPU0mb3R5CS8uxdaamGA2
Kt49xCiICPo8GWaiyk26B1+n2cLRnUmjHoPpnuyR1FhJ9X+U3zKXsmyaHGKdzQ8k2wVB4rFEDG8c
OenSy+stQL7GsqHXKZNlwFSRltuXECWN5m2iE+NNbIFZkk/gmsTqK6HfQMNzfwSWGEyA0mhQy748
6r8p95qpgo7kUiHHp9JK7WuzdBCL9deDhpVKcn97BdW9a0LMOPZQearTCXnUZwwSGjfNCOBW7WTn
sYmJ8fZBYHXBEFyal9FheNxkrBN47d9pu6HuAda60vxD8/QPI/jc9cnRmXFkp3+dZ63dxvyXDxjL
BLMwKayw27bs3CJVFDd/KWEulkNYdEq4TTzzFeeqOuh8NZo5rUHeChh5qCEQuEevjE6HoiP4Kbr6
v8+hmFh3DGbJ92jW2s4zKXtrnNMa7l4TchdssH6XFIieDVgDzFHxkHBGmSbrAM4j0JcxZAS1EVE1
kTqU++erZhLSQJmvZH0kzHdx0FM2rGC2CaCOk8YcC4l6cfDpjboJ4oOowdk0SagGimBXEqwd0dpH
yEnw3zvrOjUuqQ1Uaij/1/PvD8TBV/64Jwg86besPRVdy1F2EPkzWUaH70LGWRUCK7Ms7gMqSKuo
G/6fLTBE42Dq2/xw8jcj0jL4s/hy/8NsdXdZx36D0t7UFEWLx294eCkuYxCFMyU40mM49JcFfyC8
spF6t6xeX4IRgD4zP4zNu8sWRR/x8NSbH2/gjy57aHIalhnEe5Ob35zoVnWiKUly8XClC9wxsBcA
VQOAwM0E64IbkcxQiUHq1cp3P2LpbgK3F2dyAYtKIPPIrTV8mz/MRmNikG3RPjm/Xk88hcveltKF
FeKr+P0pfzRhMBOvucNImr8gfQsjHML048+mXua/kBJy0oibfksoGPmpUQ7zGBsfjLtSHN+XyMVZ
QIe02C5r20GSVeyrzWCdm+G4i9GymWGSkyEAfQiqYRZtSOKVgRL3J/26LVutMHkoIgMffw/veSU3
gh1srDIB8iIAL3jcH0QRJb7P7/10de9T7ECHP+4mzkqc/434Y4XeTWYZlAiVcLUCMQRxAC5AYuqM
2lF0oeoidKFfwWBn0IxVAbJEJOQIf02W1kCT43MMO7gahTj3lYkH5ArjtnqGvqjyveSmPCv1BOnK
Y8s0kDgQJKQDsXsYrJphdmizii+ZPH/7RiaCaOrpHIOZVijIqmna3mngKuwhc1BLfGwj32WmA4Jq
VPwDva5FcGtPpFM4myTelx6AhHaJ6v7iyEithUAy8H3vHLcQklFLNsrSmGlpOsok97H3cSc61VD+
EmsRNL/7D2euwHiNBYe44m30sFeTajR1tetC5PC7eudZNgZagidiyDGtP9EmJkhrfIqb3BR1enXK
G7f9S4QcrA8Laiiaxu3swOmjXYZiEJC82Fn1pZMpchsQvEiC55UlqnlyPX1SJ0h4IClAzzoeTcTL
6OyCCY9B/xhI+uu7v8lWXbQy5y8nve4b4B7QifnrXqh5xPTwjVdIdzlT/JdKTQF9VhWGfkYC1bCO
b1onf6gNXZtfW1dzKL3dt51kLhgM2P6ATv2n9GCl7T6L2pv+O6LpJeCzW6xNapV3zjpf9U9d9iYl
a9oA/yEIiLGhu8pjyPJ2w6sHW4he/2i3Aq7geSImzpHo29teUexGWR2VrLu/HZftxqNt2JWOYxV0
J2aSLxnGqiDuvMerSBJteVUFVN7k1GYhZE2tAvbcemTqkobW80HiSNCLmrjIfuflT/xdLqkDTwUv
IHNIMHZ9+yL083uz7+gMlT1+9k5e88iLNJfYhSyIxhesnvsaoNvv8OMNjScEsbyl5QKNSrZrqMsO
HIxNI5A74mqVWPWLPGgxv8WZDAnoCe6PakV5w+RqreRUA7NyFmEyM5640LQo1+51ZNp/XvMhie7I
PtJMcz0/C1twBr70U5jGIZr3H9VkH0w816r3UtyyQiKafdSadJoWvnm7iwJuVmOWaC11s0WnkMwu
MVg03wHeTALThO8EF+6evSN9b58rZP2sIFRFdmIEgA4bkkR4hnogs3UWJptzmYPvAbGJuyuGWsAq
dC+oCx3liC69fZvO09NW4ErJf4HhkFxyPIaL+Zr3xIN9J//yzb1pupWDGcDy3xAtgvkdeyE/kl3h
zLhSd3d673rdH6SmxZ3HmjauZG7eYwG77XbupQ6RxgBZzFQNHL1i219StO3ni2FTZYf5QdjdbL3W
XGcKIPsYuh4zvjqkMcr3aqE+UUWO7L6HR+4prkIjkS4t/Mzz+wKh8OId0gVFSL3Qfq+kKG4qQCd/
97WlyUd7nsIZzINjfbbeO44W+MOBcakRxEXZKiU0SvoAPSFOacpqFXOoHPBV92yPKjh6Cik1Fsq3
SqLyrN5CuukW1Xn0aEkICXf5WuXxwJOvZmG37DIt0igmD/UdYttmQYbJwy/QZWv/hKBjF9+e+Du5
FyNnoNbGINUnelWRrfQBLwx/Drks9o3fbsQutvywG0YSn6eqC8mygs58MAEFe7RDluf04RVZXqPQ
nH/v+uKNT9aMJ1QNcj/0TThgHuzrFfyvuh8wlUjcjkuJDOnZ8DVaF44/LDt9toBdu5MLryQptUT9
Re8ksafvin4zP6L9QwhZfxj7uoA5wHv8ci7cASjsFiQwcPI1ZbWyeYktN4y3qt4DcRo/d9b3OCeD
UXmOkeYkc3CqW+URIDnu8LAW7L9eSvz9/eo3qTE17eeuBG3KND3P2IwPKCIDwPMPRjbYuv/pCwuq
YXLGngqlSRbu8/06kTIgUZXtAxyTbydb7iWfKq8dFQ7Ifwra6Z2bo2RDFA3lNJ7VTlpgriRyZK2v
2FEeQct8nEdLHu0vNNCseA837VralHhexkGSmeN3buhysqlhFlSbe3Ri3uiMt4Lj0RuIp+BL4A0t
XsGeb+4CKCIzv1jUtG2O+cPgWM0/BLTP/V5MOFNxOOnMuvD4yO71y89DiKfMFfCE/Nd197DrkWpw
8Y1qUV1pH3rGvh1niYXLNWihti6H6RP8MjtntAXdRl0sDtn3BJGoOThuVv2t1iRL/QVMUcV7QY0e
DWrRQyGZWtSbBuUS4Bn58dSZhXLt+x6N1Y1F49BzJFHy8ELLpKlLZzlpbgb5sg3hGgtF8C39g4bI
Ak4AxwU1Aos8TRFw8g7tclGxgZAGrtxN1rPMudC0ucnD8YwBMinO439ahMBuFZj2UrwNqNwldNu+
TyFNHsU7Bf/4RTECENZnlCbR7fwV4+MB9t4g6LTKxbceyJ0+jrTVe40EjVYD+AQLFVKftYCQDqvU
PhDG3j5qaa0iUvuG5iCK8Yg0G5EHLLW0u+rF0MAUxnIxcoWO7/F+cNN1bD5LvACmRvoSDVlETeep
2k+2aU2f9C0NT12v1/BLP43Lwjx+LoUKYdnn7OTXTna0FMp9p4zp/krMKq2iSAuYnyWwWRYxDdpZ
4VZwdpx6tHsEx07jorleVX9q6lToo0vWh+LW83GEUH3fYYrdk06Oyg8op5WVzdjcacWAJHtULH88
bu11HezxeXLwsd1duEGUk6yDo48W1KbJiO5GmbUN4JJnCcl8EiZxwZdiLGblwo2N5vxBPk1cLr62
6Zkqbtuf0ZEdqfc1fGJBjM8g2L0kUBnGqGIYMXYW8tKQadjojX7WesrImzyhO+EWVMjT1z4/ot+b
od0ew/LJW3B/Po6OxpQYXQ//JDYniKop0vuyAvFv+obV1BDW/nSpiihZ45s20Az75HAh3muCVhrI
aAqBHB2ggmeKjKGfg2jXegLFm17I084hGnRfsn2uh4j49Ug+QIVO9b7FlusY+5N6dg8EKTUM+/Oa
7P082rwsoL80Z/JWO4afUpxyh4TlVcPkyuLdv5UikYy/NAMEgNMEEzEpcosc64pNHq4W7Lcxql3M
6IGHGrXO0fjlCAqkv8s1Oy8l1pom3tGL/wz4Ce4lnzZpWjYvdfKRI+M8qgQyB/yGXky/Gby9lqdF
zxsA3cpBYxr6r89HfEao37ZPu+LMyQNdT5/9LYA0Ou1OiqzXZJBkJsowSqbqWy0etLRGBMh4oAVb
nQntQsOjJOifauGo8p8WkoGK78HlzQEUNr80U6x8FyaT8ulEAdZvGjtddjN7x1DUoe7ZGmnB1IQu
TBg23GlmxlZoRNesWovNOrGwxWx7D89ZNuP90ZVsu1pr97azLgLpnGGHoYAE4OdxhjaP/Jjl+120
8f+vOG8LbcjIWF76fzGBUvM0gPvwMsZ3teQUhzSxtvqhAAmtA9iRQZuJ22U5XIvf25kdR5Y4C0eS
Yq7A2S1Qctxsq4BlzNzC8A6B9XeAq5xOrFZCLk4j5K6aLC7d+FtPR4OtDRWzqkhKhP8XnBEbd5GQ
MnJE7/Ya7wFibpHPZgmGCEdarGQDCc5Pljt+QlAommthuqWd+QOJV81OlARDVqi5OtiCDRxiFIE+
06TdDeKej3Gx2i4PdJV46W0kUOHqFDAALWclk5rDBSsJ/xWC/HbOXT3hsre7R5oJv/Oq/yTSG5TE
QXBMJ8ZnAmYNjNlIOR9kKuV124ApaCt4cbNweAyO2qH+IKUoio/wEyJUgtrcsFONktHRvfAJ7qXB
mCQo91DIAGb6BTY62HPiJvYqwbZ6nOdpssWdi3Wqv7fhcOD8GiFQrNsyNi37daGKw31gTDYFbsY/
o2CpjAQZmxLQEU6/8ERuoVLtx4jmF1DoTnLn0p5rbXWAvBesDtuU8Xn2q0nLJWlyuhksnObcRQCq
zP/ZMvS0bPUYBDk/RYj4drIjLs9DMGyfkD3n4iciVYIoRZFmnQSxzIcBTgcQ2xQJ6nsI+faxoloR
tG5Csr+fft7Zpw/e2T+EQZNS8eM6BLWwBVC6ClU+sNceprW8S4bIipFm1558beQtLiutP0YjahhI
MrRae2H6C0kf5bJ1iSZMpaLCb6IDtGI5sCRkAeDUZxAk10qrrzEselSViaP0S8q9SVcQEJoAyjkC
UFphMCsjgK4ip/3IaBr8WwTkUlaWM0U70oSqPkOvBXUR41W8oiy38yPW0V69xUuZ+XciwaFTBNzn
4WmhCf3/twfzkgA/Elq/ZTl8Ev0sFgjWk173saDkqEZiPUdrBHNkpUTuiRcr9OptbBp3THuYTUlX
WtibLz0TmPxRrqVH5X9D003w82YzLGeU+Rt7xeiKY4LVW1vArpgmUTzhCKAW7GxMaF0U8ybWdcLT
nQ55GhdvvjIsb0VNicAuzNG/leRd1eIxCYd1J8QARN2O+HROIZKDPCj2ARX9netk0sJgBZQfSvLh
vMM/bHVkgYZFpv9I6yVHl8uLVH5WwOoTiRam3ctq5pbXY5zjKxLyqz1Yaw0A/+6w151lvLYUk1uP
TwLJj1dd/jdtQP3t88Mz8YKFNdeHPSM3W0sVpBvgmha2dUq1cqFc5wNTCAgZVHGwruWvj+YjjQ+s
ZjQ9OhXtVr7nRZ1jSEhRcoac7Yh043O+krqVO0r9LK1r9x9dbLSJw6ogT0zwPQ0KJdk+qa51AOaC
y+iMajk3/XBTUQSxs+c9isrfwm9i1fQ8168jW9KB2O+eoyCElUeZShiK9SBGMe7lZe5MLA+iprdG
KRqucN+3vmdH2Y8khj7I9NerVQHtk1sKH1lRcYPBChKRQ6Jt+7/yD82Bm7Fb73K6fzhTpFrIB+J2
3KIWLIjKIFDlF/b1Y6KZo8HJmHObFgr07RdXY7S12uVzSELi+xbNi+RNjsObkTVykhA2BevI7jGJ
e1TqlhrWK+c/O8V9r4lG2XG6puFN9vlZ58GWMUG2dK5EEmOkbD9FT5r+kHQbnmD3NCXdkjgG/zoD
GokUUQux0CIuD8mu/rRUPYVl4/OOGUWHGzQ3n4Pal72cd/akuwaMGUB1Cm94QBVk++mRPIB0cDeO
HmxmD9GTuP+6Eb6bBg0nZJsA7GM9o3v7xvqdHZ+2uDU6vewMNFpWGEeWQU53IDWEsGk8PfpE7ZOt
DsRLWhw9TNuQPOOzzKHlyTmcRmkVkXzmXvI7L0clNoFU31ijhbhbbsrV1N4xH4AuG8HuiBbh+m4b
IwfoifIvh6lIQ5cefD3Ye8MitmW/wnRIYxPJYjJ4apOwap5a3OQM7LAFflelcdTRUjGrz/xsRXtC
fj3OC22d8cQaA0onVaIlJ9KfaVkscRLS81OWsxm+3wFj6yvjzkJRfVornjw81NqKjLYpjz7l10HG
1vpTgN62vOgZ3QdaPfiqbP+bmRSoD+COwe1THW4E2+fjIVN1vW6VocghwKnXngNzMBS731gNA4f+
WNoNHwTj7uumWwuxlElaLqJTsekQtHzgb9Zrikrmz/7NAB4x8ZQJoLldBQzOgXFBvwK/2KsPWmVc
9gijB6TvGUwnBJscUE8CvZjlAup4GSinxzJg0i11v7h2ZSXFB/2DzmT7hO29OIqAOU+Mv2Z7kyGR
DOcet3LpYPrenITlsyizFP+xlAZ2MoNdgxddkADNw6HCl1jjEPCR04CQB6PagcmlsynEZHNXf/64
ODudMxIO9D9xpOtnj/HzKHJBFa3t7c17kMPF0Zr8TTARPrQarB0QOPLPd4czaXVXBQgEoeai20AX
Mq/YW3b/doXr1oO0nYVIV83GmAa/92zacegO0mF27mft229r38nLfNoN7h2I+EtcvF+4ASx4akW5
TfAQ4jr853ADzgkKMAdw0DzzNz00otmTULzb25K7dPiUQv8gxI5BYPIqSC+B3e2lAUGwKcLeXt2u
3yi4QVXDa26isZZuqHTX3Y+6kfl2QAMsmMlD6K05Vn/MuKPOggki2HSekTPmkhHYu5cF76GXGtbj
NSf7xESRMVXoloDGprw3/fkfGHiAjxOHXkHhB/GeMjUV2dtvPyy7FqY3jtzs7kLAldkfyns6AT6N
Zj5laDC0SLay1y01I2N7mzsyq0Oer1AuH486OJMvmgh4xvROS8o/HPCpIxphx/qGCJ2tktsrlrce
pkLnaL5DJm5eylZmudQ9Ngw7888efnzz61WtbiOaocMLMYj94tHbo1o+K9nShcWNuCeWhhOI40dp
Z4xZq4h+JSiJE7osweZQc0BZcRc3oRcbtZLeQstYXS2UbMdvQ2zfVN+12yTJZVkDB0hD0fUpgEzZ
otwuBIXzfIk+PXS0UUZXLQBa8ZU72Tp5V/GyJcmyXq7cbGfxOlSLvQPNb5KtZ1omdYhQILjWYeEH
TqT6jH0vVof4MXgcQUqR/PBYC1NvVS0zxaFH7HkXMVE5OppWYrgD2cC42Sl+L95DSy5yhYQ7riq6
F4RfvivfYFPIDd3TOPaiQIiYUMvK/dS7BCTpcH0D3Q1Bj+1BSGmOisO9yVxvhl9Q2FvxsQxeTXH+
p2jeYJKiWwQaoFqRyh+8SYqC3aAdRj8nfwZVPfOCgxWcSIIO8krygar9SeMnY1vM8xiK0Xqwlf7d
bNvtwmDl+2il4RI/FpzlArIzQNmAql1GAxZBcupjMnSqYCxqFab/dC7HBmsCbInc3Yw+pvHht1Gn
qMAL9yQ261ZggKcwpJKVNiPh4+WnSHIpbhZvAwTxL/zaeCTFxR3oQx/s8H2tz9sAALsXXqQcofqh
y/nbxlevFR0xO/RvX4Cr5zEP10lMOqGE0FEHF1zBjIFBEIcLKgxiggymxnAKJBD9so8iPc8kB6fU
kuFvk1cYdadP30je/xAzzBnIA7Hr3Jz5ybInyZ+INdNkYfTzAJYfut1sJmeExIKHoQ+xUVIe4qYV
AleRGZ/ACmxxzVkt6QcPbPw1N+cV/xas1sRsmUQYRz3ElcHhO5eACft4jGvsnQ4JgAkXUiRNLQBk
UU3tIurpn5vbndNkgni4jKMpqeTqUyQqkbqoE4y6LBw7M8V/gIq4Po3r06LWDFDZ5Us+TrNIaJTc
Km8AOb9xZKDf2cdYeV+f+ncfLb2PS+NLH1hCRBsKqCFK9bojZf/Ol6UpJwsvU0ie2FiXE8T6rR6x
WsUz62whYVz76knOB7L6YaVCg74z67e6zwTcHrLsC25OFh56kW+6D68bXcA3NVgPezv5KyAthtOW
rPAifkGzNiEQ2UKqnQYQDjZTdsaPAwWo4aY1H+kIv4MfUfVGnAqadcS8zxoQ9+qdJEzQ+8DJpWhb
gD/BhGTJEK4JPQPq4pHGXKi2x/gQF8yU77vG8FMt4GRD3QL1xBklSZu95RcEOaVPXCJbipWAu9e3
eP3MGQIdwYghWAAPuG+sgs0kjv283vkaRxkvq0Q/Xg/uI45Yw5av5C9IJyDI07zh9IEqWeG2Zyx0
6gvzRCQqxkZLbciJ3u3xfLMOIHOBs/8/veFYW3CGXSgGzQW5i99s0VvDJb6M7YTv1mqjHPxAqBlH
danKCukY0DDaZ3gnq/CoPmuZK7+2VrTHK5O3jiEmh/vy/0jK/Da/4K7tT+blUDsa4gZyiFuwOwZA
XDYjYFj7etSYo7PCyD+2c2gDk/C2SK1AyFKFXc1OKwVGsXSWWapeNuYKlejA64gn510H9VaHRD7D
Ns4ez3Ouoj+aEVrJhI9oGSctpxjHg+GwoDEB169HfYWpq0mvLOvXG5jS80WoaJdnBTDImKiUcdSA
eDY33ahbMWpz/7thKvyiv3GVu44ZMJMkcO60uf8SyrsTdeDvtImJgAcY7+MXYwtGj1B57NEjLB3b
Wj7FfADG0+d8szglSKeYy7rwzip6+oeSFRMMZmx/tcmodUquQBVWT1F0AovO2NeOSbjheAY+3s+7
/FI6CFPMICF1Ez61smtkhLc1kDESslfTgcETc9nZSQ2Qxa8BF/oQAAxCAutC1cJ6yHvE6i34zKvX
dpAUKG4B0nIXX1T8pbLnmAbOB+9ObZol30bp75CnLHpOc3gRbPqcXSIvrmQQp83xjm902PYJz/YY
8RqsM/y7tewJDLL3EbIClHR7dHecks35GsFvxP3bAyfohiCHW+FQakDHgQWUBiIkowdkP1xaI3em
Fd+N4P9npqM2lngQSIyVvwwvdDovA8/gwHvX+Vyw7eYqsAejefvqTUpg6urPaAy6tUhJCINr0xEM
Vo4yeuKd1vrvC0nun9OwJ9WpGD5ddodZKe0AyUQu5F4aV+TFIqrqlAxHKyQasxhCFGz0DPttG7BO
gpPqyzsnC1C9a2iS6T7+gZjcV9hojxvPIrj65dexzJIFZ2XQIYqkXjvNxp67mZjcyJwmOst7aSUw
WW6UNdlhsqCL/PWQopUgpr9mGV2YUIzpQeys8Bc3DxfmF8lolWxXRzoQR7WA21yBIgiEU7n3Egwv
obDB5+ZlOucaue7/JrRpajjGJpfEs51nO3yD1KSxoWLx5pWE1/4ykEzg3f7ZrBEUMzhKCZq7Tk7E
WBA76or/AwfCZM+DMwO5wfgTItk/QsH71M7HaWrSNFKIAiRAA5cjRPEiUZtyf/VXx4K8lTnSHkur
o26wHSkqqdE0pcsti4qACUcFiIIBaLhDNGPj9WLAgD6CAsd0dXJ0t5+QQN4DDPa7MBG4UhWZ/OzB
+v841TwbPMLHGCiCEikD69n9p46cx/m5G8Cv5P2SeL8KURBk1FxCYc8h2XAfRiwli43FPX4SfQ+7
6V5AY6BS7OSFd9V+S00gpYjZG0/z9+KLI9VQTpQwu/yFKoRcGe++9c6VcL89j/T4DJXQ5grbtRup
C3XYQMVsoCkurOxFyPgbiqQJGUsME3wdAjQsezpZM0ChPEXnmxXdsYXekn6fvjD9j0+z4529eHoe
aXVFKY2b8ju5PHSrVw7QbFPPnQIbabJRXfwdDwnkeJHwgzcXqoZV5AGxUAJVRP8UEq5X1jcNRujD
VSs1BbJ4+UpdQz6eeMKe5r981fXUlZ6dpuvhS6mhnRsElv1Dcl5JgSULk8CCfqjomwYvOSwTcrJR
gI8XyO2yvpV/suJN2etlr83WBTKuHTQYqcs1/zIdG/wxlz6n7y/w9/tLmHnf5fsEGvqgDanDWHnO
jAMMypxQ3h7i3rAgnGCa5OmOR1zTCdqyk5oOcuCKVazBAukW4xw8KR+A69oGHsERD8H0JqDC0vMS
KcMypVvqGxoqgaTfhvUhaMyptDwLsGMh22Y4up+QxLKwpYIWluc3hX90etoktSxwvZPL/Wm/T/Lu
xHIVt5llJWizO6SK/fmB9kZ9N4OS5lRoCy/1k8fmBZRk70sRMB4bj8Pi7P0XPHmDe0a3gBcks1d6
V3gZoxkd0toKMlNmBfA//y5er8b4ujurd/CyeRi8OzEmvsioiHGenVxHyvfnCObfIcIl+oQtVkRv
Wz2fr+BvSc1lTMLZ03fa2mAZmVc3Er/Z/ts7Cx8+gb2hlDUMnHau7+YRnRfp4vER7q1j8zCxJzGZ
mZlbXgmrQ6SND27W0E9hSFIzT/zMe1yJWUrGYyGi7nYspHht86OjXKr8ZSWYzUPklj2MXJTUYbcH
E0DIrW/IrZ2k9RvFIKIzCJUhUjcY3iH2O7shdqkxG63hj5NSIjS1oz6Ubi0GHfm3TleRZnIQdogd
gz6mkWaB2lg1PvwymD5CU9VvCOrMYi3dpDn/d1wvzWRi4j3ZkYMy2PGb5Q21vRJfSB4Q6WLrIk7C
ndSL0gegyWW47WmjDaG/L6z0jKdWLv+th8KiKRGAr3lsi3EIzTEk1P6HhaQjhXGFFxhMiIf0ybuB
zuVvomLbiq6AkQ9h42Jlc8hW5U+F+k+eXPj7BGrci3EjikE+aFlbAbtQQ4KRZgb7L5S9h+pI2VdX
LtYc/zjAJhVNaeV6GB+XkBJ7DLGS/4abHWio6MgtPrKe4Wt498zCahPUBb6AUYcRK7Pv31F1ZndE
WTTwAWXRlxoasZhq3Zs8TFfrICJF3zXxxXtkhT2WIXDwZBSQ9Hm15EwtYpZvoeaAaAwFQo07fXE/
pDIuPe7xF7kXh/zlPa7Wz1ZaYF7CehR/TIn9G70E3hjv/QmH6e1ZTdssun1IiBBEueSI4XQRSeyb
HorAeKVbkN3EMdD/hqLpZ7p5OVoINo+B6/9Fjym5ZxM+jI1qPus0yhBD4QKJ8i/jX4EvVBtavOGW
09+qjCKRXbUMgn6bwh4k8pFWS5SJaxekmpjva/cEjBBXvVs0LyxWoQmYtXhnueAcvezyAc3JJbNS
WQoIN0QIOs4x+YTeLaHa7UWIrX6Mc8i1haMMhfqvunx9RZjiKfxbVvd7o8ct9M1XoaCWOejtUmLL
FRJaFqLXa4HdESDts04RQTFSR6CHBGbuWim/tgnOOuIRcg9u3ERL/NsWTYkYE0HpY6/8i+y84nDI
1bdT5BnrR9/lxrsXj5LJUUlK4D1VmBn4eMN801hvW56jSZ437GhlRFcmI2fQo1I0T00THabEJyJf
LsMlDy5EZwB0f+zKNmfSehK4ETmp3xUyoqvH8MxkdAbrB3FHIfPlvI6Ioln/zshphVbHWOtJ2jlL
L79bbyus7Y1YGALEfz02gOvgKbvoqpvWAanzBpGpL+p8MII8Rkk8XFOkHcEFGHBQEYgqcPF0a/Y1
w51jOnt5vEbXMDqrsQ9fhs1FaH2NNcFQ4REQe7GvdcWAoHsU/lTpr8++18T0JqXEfZyR+t3tueLy
eEcAilyeAh62H7kUpdUKP4hkNN47DrFalFB0XsUThu9LcY6uoHbfX4/uEudOYFMnlSW24x14rMwp
9NpvrvDh78cfcCTzRx9jfnu4Kfg317+m9GKUfOhXtbITbTvu8qVq/PHdubEKGK7Hve9E91fD8b7Y
abQAPJLopijWHu7SlMc0Poq3JxpQOvtN95OZBMmQXEfVnuv28owcJJgaDQQgKuRjLvj+vyn3Ge6D
E0rZByAmmZpgqEh9XJB9bs20jhcm88Ix/QCMd7Mb4E0N/iWM3yRWaYU1o9Pfh1MpU96v7rmeZR1E
mJG6JJL9LITAnFYtDGnSTFtxiB/yN6VQntDxYNQtzNBJCU3TdTc8r04BHpGkBG3suOYG4NsHWe/z
W+URXcmIdgXy5aNYZRDeZeVNKWTXnI1SZNPy+yHUGDOim1H+51xZnl2yB1lswXTNOGAK0PsX9sA8
5TQ+qB9wWIc6YWG+beBavcGm5c9zGYYb+S0QMrymgOw3xWeZmlpj/JjoHxK+LgjEeP2ctHr4vykb
2iALJttsf2/3H4jecW5taOBVBdBz1Tg87yTaORDtB9Jy62T3YbksK/5crlA06XITXzYl+WULgLwj
v/fi0CnJEnR/oaDLkhIY1H+CUb+Yz6UjjSVLV3aqbLXoKHITymD+OJ+WHuoTpkyvHJYq+sWqkRlD
WAjbPCr1c+EpK7ThsRNmGToxgAVIQ4u1wm1QH1HsDu9dFuxT1vwTs3RSM5M621SYUegE6ZUb+cT1
OOMU5eovjyDXqqTPjvrGxqIYrgYoaRnl9eJT3h8udpiTBSeb9yQNcOR17/TEmgPXLZQUcFtr3kws
Lw3mYIXhPavzBk5nvfnsZ4TGbcpLxqZOpDLwoTM23mT5VCY6U6m4FceUQ6P+TKKf+yCpGNKE3CK3
zuwV/6s0GF3WaRT6Sb19J4tSPaemMxg31rqWGtv32nFLWZpPCaao52Q3vpN87SGBLaACEEzFTdpx
UcnTddIrl6Mg24hSV2+PED7SauyRR7PBkav9oJfHsDOn6AzzARvgSTjSLZ4nP6AGD+J2NPyAittg
+H+zZmPkBhgUQ5LRztmCBq5nRwBDLdO0R/qI+dq7c7nQqhJRM/RuvKb0d1JTy+Scbv40e2jCx45h
4sNnG2wy3eujM8EY4fOweQV+P4F804BcJKmG639p+LjAdibahnmHfx6ukTI/81JFu55QbJrF1O+Z
PVRYbRPXVOxbBnILsJLg16rNcMgnTvJtwsq1s7SuovHd3F51n25MuTsPxqjRH2g9u98xvQ5G22qs
xsZuEGwp8wAq3d4ay5fEzn9Rpd9p4XyV0Aivg4naY/NQrDCWYpg4lggdD032ihudzwIMIsN6+MdQ
crTUhdXtDJM6oLnc9GuznDEb2GWDBNslrVZViV4OwuuWVcHuE8Ee/iSlwj8j7LFv0EkNkFsb1jiN
2Q7y+GBSHFh9FYwUZ97u+jOO74nnFytp8uur1RAff6FFK1rKOpXiFOHL14HEyt0fO0CeP9mB4nda
xQjSOMvreL0zM7GGHB+85t/LmN02Tt0NDJp5+DUbyxI/DZd7dKKfdCmYLdeQfnxvOYpxJnropHBb
6EX8cZ5KT4VFYNiRtmdMVWahNZHxOzItMPW1sUvAGXJ8fw8BvrbmsBPqFw43UqrwTMEdQmdWc7Y3
4E1YEYcjEc9OuZwGhGsa7xtc2rSc4yDWKdw+BEwtk5QAMTez51MOkBO3JkOOlL7zJcdDrGij363e
lRfidotfoWOrdvM3FuTPf2GNEusOXaRQ8Jnwpxre3zp32lv0+CU+lanxWMVYO3BOZNM3S+51CDzh
AcI7l9eHV+Sm3rG9fOzvZirmwpY9ZAC8/Sr9S7JpVEBfrktTWCW0+LFpPT/a3I0d4D/eGo7PD5ce
aOnW0IiENJ0U3zsgVHZP2I++vIrcVADv5k/Kp6pgqV0C8e2mlHKdv2ZPF0Wf6AjmDFk8oH//qiMT
Hhwa7CaeQLlTSyxJvsnDdpMHHN209Y7l7+QEVKcBMgLsvny7jyGvNgfxlSBe7+IKwAWO2HL37XaE
1/etLsvrfQ5Bl/AAjgmAXcFdxOoIyHcxEFPWflLRB61XbXDluNg03/GslNldl0C+xk3NtATfmiWf
DiV6GpzSdoEq7PnDY6cpJYbYzyMJ5JO9XNSqjlipUCc4OZne9gsPWVIxCuXOO4ckZGD0tPK/r10r
7NLjL1A4ZzQdhx6rpBS+Icejvjj5CB9E7ybk8B0FrVjbfSR3gHcE0IK/mrXolTyvsJ0ojpfAwoVy
eWOICbcY2PhvwityQyCCamkTmMcIYmj/pcH2ad0wpsvWuKOPnBeSXPuhNrXKSv83+rm8fdGSd9dB
tjTuDITKXFuJpDRcgl3f05rSQPRN1+FJWQIRHbYZEBDY3+tx4zzsdYXO4typhEtaBl1+7OiNna7G
4aXqy39BZyaiGXHMOCLQHFiPCe6kUuLGFnLvbt16tEqn8kvIa04kC45rG03/5CAtHJOwJHcH9CXx
keKlLXF7UOA35XcpqlxZCXW/orxZjBgYseoiESiC7LHSwGVAXDWevLCSJcdi8JSa4n1/yEvX6NRo
5mVaN6FoGYhbL5NULQ4djiHFSep0u8hYJeYk4aF1Mbsbnck+pu7GIzoALfNfByWJFh0sHVfe2crq
UacSy0VseRRWcdx3B3mLVOkifE4TOc1VM15sL3Uai9ehJXzUMDz3t8PNW4JKggMV38bR7MI7Uedd
WNrpfB+6TDibiuDcNv8S7qxKf3I/WsTki1aFyr/0ttJY2AnNw+T8U43TVXLTEttgAIyRf0n1KYsZ
R/Qw6mW0u2Rdbo655zNMcknfyu7GcSEeI+ufyu+lIEbb8Wke2DEJxakBPtv2MzScqKLuPWWcxbzB
7Q/JS2MXAmLvLgGdfMtoufUCibIil8r4ZIl51ij1q8KSRJZ4ahxhxOFOENxSpFj2Hv5SPZc6+Q+W
ah2VVOYlqxXI7pw1cVhjOdF26XmH16GQBRBG0Wo5c9jJLaiiBPZ/6InF+46kuBjUFtMQ+8F8gYB5
Pw6py1qib1e8cQ+85OkKOjjU+9If6CPpaJYF373Yes//d69T+f5fsS5qL7wV9tsxOFH+DqCTWhUc
fVKDKc0KiDW5ycruovulJgDJ1ajk67LZ77c5EIM87bQSfAj4hFflNAo9cI9J1J+kAHrsVWG1lEXA
EOBQAz7W+PuBopzljIN0Qb59go41SsEQqacvYt6rPC3w/bgpKrC2CQ5j4mFpAb6br39Ns0NCq1IX
xxGtPFAnAcZ+IDrxK1Azl1BL/W4HIc/sXYRjckGBVW7KBf2spI2Lb26oaWbaFc3kpwf9k9rBcTWZ
J1E6ubAKA79ZtU9UI7KlWnjfAZWwh61eSfEzoOs6RQcgO7j1lYq5OWzg4z0uDpfmLKAbSfzENbYh
RKsJq8pvCZ5eui/xzOeA8GydrZPjMKxffYtjUFpb52W44E/HsN+/V7hVTpCVVT7bi2MAPIe6c9Wv
6zMcSDoJIMvPs7AiD5UudQKgG4DTdQeJKRdX+bFsvcda8KzoNbIZLrnWFUDBLppZVKx+Co4pJM5o
kSC36sxb71BVUEa9/p8xFASLVHitUrM9tHDgvf3rdEF+0mudPIcdrGyY7Ebloqy2DJL3u0Dr7xYh
1IpFseYChEPNMrUOxpglOrJeenh+p3v8lpQzFrmV/lon6ktuaIE3hDk4Xeq2BNVREErksJ/m/VUG
Ok/39HlJZ3N4PCVzMVn5RP963MIfJ7r3f9jd68V1UvmcFrxjjaDBWQM1Fg7y7uLQKpBjAiAOf7yP
QqY+sqAh2Su1W1yr1qLNa9s0VU9HAo0IejstF6etl7RJyBxRRfyLLGOfRv+Yfe1PJkqj9ETXj9WH
3iXr7V2EUFkc/lWq5RLKGrLoQP9nD+C56k/RfwuyBaCV+xWAnlArpZOygQV/Lxg26nQaGv23NU3N
6BOvye3N6QBCQLUimUPM6TRmfEJx/iXTzobHNB0c23Gwbc6LYS2dsVltmKvFO7HEYqqqp8vJRVVK
Xevp9k1ywTx/9BPD91vjYguGQQFcsm0al+52bsWO5+Mrq82OLgqbMEOmTNnUmkWDrOu2bE19aq87
WWPvdw9IvPOxu4rDtLO91PkDIOMS/LNrz+pRuNoTI23pL0O4xJm+TqckGuBtSYTCA/DvX4Gw+JAC
MyagLWTln79p66jtwfoepdjuN/FC+uCYkwKlL1I6VQU518N2L01tmLJCcdcc6VWKzBvdbZhBskC7
Xx6Xe7lI6/YbWNjLTkRjLlvhT2at+IidmwlxGV43YvhLgXhtvORg8f1w2hfV4MgxJAwkSd5YHmoN
7l1feou+peL34gXHHQlirV66pDqmLNb/HtdOSZZkkL9wWqflxyHuNP5fVyvuMRJ2PPizYZxWb5Mg
PO17i4QntNbfWqJpOnb/vIv0I8hv9+xIaVOVfFhnvMN330b0KD3llUhFBxPDj+vJqpNp2IPfn+jg
wFatKAmrDaYHcLISWtisJKA6pc1I7uG4+BNDqqyrH64xxtxvPbNBxgXPGckoWX3hPEyVjqsVlcum
b16stotx/c0yel/JmOSQ3mWZTeMOe1CYa99/cbT7kY2oecFiZEjhlD0XXb174jEW/ow9oR4d3snR
OSHIJiBEthSZBoOxaVZIbctnhxu8ahJA6BY3wdlRwZiDQJ4ZSt4T5zbJcBeT7rrFKVWfbSNSDfnU
IEhi5/NBU3BK2Z8l8WnIULmwipDUWIQoHDMX5/ASw0Ry3ldkmyXwF1rdq4Z1g8o4qMkh5VEzz8Rw
6WmIFjzwL2/eD0uWKUB9kmQxCgUDSujJ1W5PFNwJRS/QoDFTlRt5lz9Xdg3rMFlLZrVRVC1A7s2i
GD10uk8mFCq6TFPUBQ4bkbzqgPVamvmwxIFzxYj3EMcMyCwVJkvVKzd5jTMM+QgUTRkAjv7ggqro
sfu7pbHEgHICaHT5WcQ0LJ92PM5n5O0BkYoSKYRUWslbmJx4ns0Guxy1z9pr/t1S5gOufd4xRDu7
OeLZan3fYMCVQGveQXsQGJ0ICET2fSIPkCtzbx2232RlRqZTQwrl6owznl9iVMNPstTWreF0ts9a
/k2YiX1aLYPNHETWDV42To3VwqKpjxS10+52NOidRL/h41OBqp3rE69fH95GSiDy/Dsg+UQlovw6
AYtNqjmaXqEV9wVdic7+VsW6K5qKpJu4Jzf1G8fseeIkVF6CBIAjGzuZIznYvkijNmH3dDKxbykP
J19l9Vj4gtvV0cGNMf/h80LwzfMTCXsAHl10TzujzoEELlGSD0+K8sCDYPhjeEfaaRq51wRhIkDi
4LQLkppOYo/caUica8QzhIjo4F4f/z4FpITIq8HT2LFsKR9uyKyN69yxcBRjg8u4r2TOYmJbsSle
36GAf6Wahbc8qW1Amf4uUpClGR0eIASrGzsLP/0nSJCsLTaZSswcBV+CxnezGsoxSG5njxlyJ3d0
yf/xJNHgsvYZ4s5jKZ4cSMPLmt97r2yMa9inLQyS9I6MmZfd4lcs5qdU4qIiehCIxs8S64DgAaNT
kSfPjDMMJPqYBAq3DE38vyNbK10tDT0MkET0rsapaOZvWWODipHYArFQRuMauGH5VcGx8auYs2y9
iGeIF+zjferFsmniivmzatqU/7m0yVMikWutbykiKVrexRek9s/a3qji9Z7m/Ft67nnWU2a+EPgr
AgqIKB9ktYE06LJTvMonR8vIAxZq88g1lThmcOO/OHZIcPfMnzaQ3RiJpG8wG5dnL8mRohyWvvA4
lyYDrCvTCogCIfWcshZSMZg1PQsx0N/PnI/PL3R93OwdQke7mOL3D7rb4P5Lm6vqx0/YwUCIVxA0
Lox3cDH4rlVqYpmvNTmV/7xKxmbaEBe5jBItY8KQIKZ62cfXAWlMgJl3/GR6ZJLiWUQNiYCUgT7d
+/pdVHaEOg9VoxN5GIlDHkwIedO6L+Y318y5u0MCLKFdq6AF19UEjseX+33UAFvTMInjCB0ZDRDf
xT97/gl4XNEj8A0J74InDHrjBPbtrU6KuDUrqVtkbqYGJrVp9qNmlw7GspDqgf+rnmYj247s1cWl
3YKrbqvzwJbsWkswi9bhiu18CFt0LDA0AQrAPCcI49Z45mdV9ahiGSIgTBVfS9ns9Rv0kKPRElfG
9pWT8DYb4a4UQIA4YHXllq/oPAocy+CZYDLmtQoFdY8yOgmwPzqS41L0yRunF76YwS4Ir7YmuYdr
j/HDKkzy5CyQqNdIB5X0sVjqET2Y94uL+jJNJxa/wL9np4V/VuUxCg5gkZByIVRm+8jOuyLY84bK
rVNWiMaS5hVXzgsxLKnLndi6qC3fwg54pNiTnMDsVFBExjPv3RYKuj251vRO87IaT7teqQ6Sf/2r
q8Y0zKJm/W3q6cbEGveNbNpcODcaySBT8av3q8LgO0yUOn0ZtwGpVUkFs0My2fd7fQUxkFsqTklD
l2b6ULKXRJN37fr29gbzKt8pzYd3h/UBCs7f+iGe6Sc3JdInHwZRtBmfmfVU6tEtpQC8x2E9QrN/
0qHL4A/ESpLxEUtiy8QVmgBCGkkYwe7hd040wLet/nWAfJQiFXvRIqaEtihwRPaR79c4XqvYz9vm
AgmcOhl5R8y4El8hqMlMDxaN2wabOO/6F0+vyHeRV5KOktyQ8HPEeCm3n+TG2Tv8duvksl2K+MAh
RIqPom6XOcGP5x1RzKEJ6HQA3k0SxWgRIoVMtcBjiNtTR+Bi+k091vc1mWVthh5RNkyml35oA9RE
SrLk4e3GqSwXErQDR0olq0EV8xneVe2gv3RvDy2CsDkd5Pvd+SbgREO8RmWL1r6ZIv6lUnixxi6D
g14ZXL/bNI7/uN5xBTiVrl09SEzgXLds03aI4w3nixDZ9D6XRQNob2JY3C7LxPqo+vqQqNkL9DuR
Pb6cFvTrqFbMr7c9eL5aOMU0FqGObvfNP05z6XR5TuruyhOyy/iLtGRrKrs/dxlRlRVBpnss//T7
kYQJDeYUAzWxGtyem3p7vDFeV/Yo04ZhdFJR9FyaenliuxIM+FPbGMetRHK1RrGsCj844El8+ZZZ
S0EC9esDI7tfa14vhb16+13d49my5/QaHcwiNw0Wdf8CalGGwf1g4EkpcQ2K2Q2ioHbu/j7wHq9u
LhdxI/9eoUvOhlZlX5rT3QIYTo+7JT+IDEzfvxhukjP5jMRGRkmY6bV2ON2ys/jYUQoM+hq7sKSS
I2iGwvEUYMA0818oEErX6KSz+qFmLW2p7ejh3+tDK/KxBNw+q/mOQNrW9R0lPmUIbClSmbxCfb4x
g+nuZpY8ZiC3PxFjxsSfr79fwjdmhMhAIiZls6hAidmcEiF18WKOwWzFCEGTXv1LACecQn+PJAl5
Fh0LXR0QG0fFJLFmY7+WnMw2wjfhS4Qxx0wcUPfVOuN0iCKlr1mUjyDGEvT5SRqHuiiSOqU9us5x
DqXkZPJQNcub3r4djCUvXycZ7NYASOCSK0okcoC+N9nnHno4c77OED8fO/Cpeu+B6LERKegwWPcM
e7oOCBuTKdYEe9MZ3ToM8BYWg4tln5v+toZlB9UnbZqZjNvaMYBaGa+vayqfLQVDLRJY6jpClmH3
EVZ1+gwTYQEQJpuxt5VmL/9iXt/jRS1iLgAj3bQxrSGyBjCAplNGgd9U5Atat3FsseQb4HyvH6AT
l3G+u7Sy01VWlqabW9+Alq30shJt4BfV9H8tPGdF8sMwss2M+S4iaEfq5FTIIroQBjSV1h6Zfxfi
Po1jHQsqTIPQ+DUOtjD626jQZvYWIDA2DzPkT6xIPqb9ihvRN3OYUvHJ+cNWZ07DB9p6aIGDvzLp
0VSq/hhkfjNOoz3joXv89lM9KjVx/Io1H7UUgOYtgahrvGINkYOLybL7hxFOZATpHnBaAY8rT+tp
prPGaxiTwVawyi1McKscWzCtwQQGS9wZiFMFxGNrYkHiWRySVGB6P1Di/HgGOD1ltMGzBMhVLjOr
2MsM+O4BGD8HnajbPcxwZB0gC6ZHIr2Mc1qtrOXBlb9lmwYmoRfT/pkoYwymI5JMYlEDlEZikx6j
Bkj3gcW+n8AYJ+EAsu1N16vKuKHr9f93Ke9nJiZ1X9vKCZYk3Fns+W2tgX7cp88N1YNoR6BjtnJ7
QLPm/A/n7ccqIYEWdLwR9HHZVSC0vYgrWL3AS2RUaLebSMGtk3h3tWCIq+uZhk/trmvblo79k/pj
w+WgI62MjB4htFwsofIaXxVVJeRfvLdgH63HOc4PhqilA+UpMs0LMlCzbA4SJUQQ1z3eZZhRNgNd
8CnjRJjU3f0xIci+SdbtYbtn3LvYfL5Bv034xNXjpFeFQ1Wrt1oLOZ0qTxgvt6W6m6SUqQup6XqH
67eHgfMitMqMt01IOGknd42RfCSGkbkRuZUmOxmlJNMDXlcIbrj+KOnXN4WxGgc0eQcLgtYzoXtj
rXxXmu0i7SmwEDyRuJCyYrbRKgoKS7+CLce3iCgLfOd7qpT4u65vF5OH1E0sgC/KH8Z31j7c7B0E
ovkLXsUggqISOJyxML5d2OeKHU90bMCcwS5kHE8a613F7ZlcYDP7AJk4avpSwcPT8ESeCGlAy5n7
6tfGSfioMKtpoi+Jbs4jt+WdHUk0mUVx1mq0vpEn+JwIgL+AsETx/EauoQbJbAGxqBa1eAoTvPtL
axUAayztEfSh29NEwJnxTC0hID7hhNkC2nrxeYoX89UZlQYhZ5y7VXEE8AyQ8L2iWV9/eCsexm3h
oBWcEuLcEEKElQyM+pDFqV30+VdT6CLl8dxfAO6YlMTuNaUru3Dc9O3AE/cm4R3IKyqCL4xbmDPe
bJWCN40zv0LzTvBUsxxyIF5hwytOylZuwaNMe4R48JtDQndJaHKC76eXeUqsphutvt4UDVGVH004
ShGqLo7EM7KdXsJxrwcdws8/AMg8mL73dFwsMtu3KEHYM4MjwFCM20f6irnPmWjDeH8OQ5eZQmqY
U8zW5OubOl0gC0gVCALeTqVu65jqtV1vbiHxXkGGnOIWc/xEP6EbLA5dBs23UxCxfeQ6j5xiwJhN
H9DsxK8kI8ONT0o3sszqO2Xh7b0FkkgiBUkMpk7dcoVAHWrjoGOFZRekop333agwMcNe/KU2KG9G
dNMk5wapBfVOoB2Vw9cX/Gp/gkldHxqIQum6L8iVB1rTMU2Xsd0F+DyGz3F2IOfyq3hTFlPVHP5Q
vsX7GAMN1fhZkNhhP+gMBWzw+90nGBOzHIAjcur7VceT0mjbcokgj1qs4Xrl6YHpPmr55YQNPco7
5fmpMkobU0o3DFU86Pb1kn35w1hptro1FEmjW3riTm0X1ed5WLLp+UOxCquykY+oZt45nq/lSvy/
DEOVhQ7xWoceyoXIQtKk4LNGf46dTEg7OsikWDFyZyqvDSgQWOBI2mp2rclZ100iAtBGeGTp1a6T
Q5UnAGbbnzsEE6FjbYtiDo2zVuDY88D662n670w0ZHADumNAlqwjZl5+jwJJsnl89AsydpY7zdmd
GkeTJoSTUBfa3T/NRkXtQyW8mOBjbcFTn+Xamwhlj+oSQwqvrRw6l2orFNWX5wa5qzYTiAo0KySr
imLeYwMNlLUwYUie6bkt9Cuxtv2LY5neqEWjr4BHyKFYG8pw0HdKYMW99s8Ta5PKDBXcUtCL3822
VIKewuHJ5MsNdq9fprz129mLW8MF7/gHYcGhz7ZW715K0Cyg1aNhIryLapkaYSd1KFfqQADiRe1p
nY0/iLTDkeAlJs5pMqhgRo9aHGVNTqQ5fgTj83xyI0uV/5ngfb/ZQgx7bfGkYJcV2LZRa0VXRwe3
q8vACwvdcBerK3vIrgEul8kgzki3nZB1E2lfDWSDLDSuYmlPnspGFNkL3Jv/abazcr+loU4jCEJW
tL0HMwVcBSJOUGWNN1pHgVSATWQV4dQD/7AIu3q9P1MgyN+NqVmTNDc7UKf/cGK1oFUE9RBIIIkp
gJnow4XHaGOb4davDllqBrLW7JYWt7EcWi5EVKNeR04cagali9pIKZpAgzTDPEHfOe4nWawldxUB
CRKJsk8Xz/pE/tnO59miYCZ6Q2m3AX1WsbbedFrBaRZf3xAyX6xx8Oi9R9ScZXe9pZ/GW+G/CwTU
XZISHKbTRsu/eIE8DiTPcKuEfBev1878pi1yVmkoD04CP5y5eREOb1t7JDNZHFtI1sDRc1x9ge9A
Bpi1zJE4hdfnP2vLlV45/8PBVIO8HKO0OtKRnBEZuRzRLEoVafaFHnIMm7pResgAfDljg5iYW8iF
7CBnAfyJ48BYByOCn6CNyqewiRtxvT+xVON4yckUNiD+KHXulEkrWvgbVUHI+FMCm6j7YggeKg6X
AeskC8OOojywG45dys2gHsoNp22mg6i7+84E8LdzwHVrU+RpU/QHfb0r5tx+s2Aj1rWRrMW7J0Li
Lol2gBkm0T8Gwb4Njg/V/LhDyZiGQBoKyu22jbZoyZDbF5N7wStmqku/sX8+w1dplgHteagLIdsA
llfLM54D54StBYhQpWikuTTavZLggvz/c9XA5pMORFw1sJ3zt2cB3ubiCnI1aNzSeRniBTHRIa4b
VzKZIG6gUZXSBdIGqjuQ095VrO7qP6F4GM9pHJeFowUVpcpFTJsoRWvWgJp1WgIi+hwso94RfC7C
O9Dfq1bX59kxqG4BZmE3IY6R6GgPRsicVeo4Tkam5AewMiWP+eMpmkkc1j2OGVGXzOduL8tFJwYv
FwFHKaiOc2Mw/UyUAy/kQgSEmGiD1mafOy7G6Le+AV3w41rDLVvDpreuhSvANpChjYRxoi8PpTHb
Ybubkow0Ln/Qjgt81Td9+CykpiZ6fFKveremCz71Di2GTHwvJLBYEd/tE0HEuuHMPSHLa4FP52qj
OscTBENsMjBqNH7bPa4PO0XquRTbNAEaAjoODa2mWHfJ4VH4EDB8Yy8lIERQ5CgePIo/fdyECMqw
1D3j59UZxNYIcdP76u98tWj0A3s4yPBVA8QiWnT2G2AP/FcUHWUt7lqkY4N4YyhFwgs343Ja7KWq
s5Bpdx1/QAbGtTvmJbkJJx5E+BWyCQwcRXtEJ8QnjjL1XC2QV+nXK3XYUzOqvibK9iXUlLHUtVWa
NdEykY8IRWVUbcWvpT5IUJeaUS014ZR9eQdEFuN9XPNhl4rtmXjUAuytPNZcR+98SceBkB7pG6qZ
nZBnDjisQl+0Luqpe+gO2bTkn9Vwnkz5EfK53lFRTupt4b/MoxVCsnYOUktwpP5wLiefNXZnsfD5
yAR+v5CQ9+8Da+PmbIgkgS8AYNHIGfWEkpsQtYwHmy1XqFe3uL6tjKvHNe0jrAVHAGTIemtUUYNo
HG+UnTcNR3mlFGWUVeL+3yj1aKZRzw54KpjLohZqUmatkvr+Y59XXiS1zl9y06DNW/Zko02tZ4+x
rUjigWikpfyKEpJeIEGFZOphZneT/GpX6I+mn1ARl9A+2VLlQUpJlaTSBWa41TvoDDgDrxXmuc/z
Q44iw+ZynCCRiplKdkgexUWhBTFPPkLZqfLTv+V6vY+S7iUXoXmmhTqyv0p+RxE66uPRk9B0xlZ5
OjLrAPseeHVjaeqBO3/zqMMM3sHmPzFKZwd0XoX+djPRQ8i2oB+kU1x68JAlueXGEY+wJ7+lbCII
sB9FFXBQL87E3RgGl2+s4H2aK6TnZPZXMRkI0hmAsCu4CVV6YiV1nk02k81/uIghSzOmqG7srqwx
dcRoAMfNsiHSqzRYq9aJmiszyKB3af/TYbM74ouK/s7523geQOv3cX3yBJ+3Ki86JVFOe8+aTkEn
OhE/fYvmpOkRwVbyUofyDpNzL8LnQyLzQyz3mR0T6KvPlghVwF+U4Hq0UgIHQBMv4K8LCKWu/HAJ
xI1QYGcu4JkoGfMRRXW6g8eVQ9pCGPxVUEh8TF3Qvqo99bwNo6U8KzMDXRRNa/KW32EtnQonVwcL
RP1KOCKkPSEoSlxBsV0kIaBF8Txy6IL8GEdkeGGYN9SBZP0hWgLv9QIptDKByRA4mCOw5pescNn+
DR+PX8lcbpsopq93zHcanZEw0p8CelaCa3J6WGA+NnNnxtjoEZcCzW3ZaIQA9m0gD5Afmb5rBce3
IvYb7iFikbULKUVEuDHMfKSWgUw41kHoAQF5f6XmptBxIb3xdkmCyGxqoMcMy374gId68xzM+ODC
c/Mce4uCj4VVu+zGEuRkwiF7mka6IOAIljxfh44Kr0DNUGgSzPdFvjtJUIbxebuf8Ch1rMof23ig
7saYDtf0LPcOVWBzspd/vNzGXxUvAxt6AA2gMR7WMmfS1IWC+DrFGPoANE9LF7RMsAoUmVVBUeAk
8qr1+I3iPjb9yD4PrGC2TnfZxk8T2I6V9+ECovA7g0IjvGP8yHK13Los5at8US2FVJvsDPVWJzj+
nGm+dTeIyk0nrEeoF5Jh8MtnA8L5AWOIr5gn5jji9HIl1NhuzLjlKHdSComSA2oWo4Sicd2Yb9rF
uoRn+XdoNDaozkwm6q1q/DWrbXA3pRtaLEpoJYVWd9mRq6efj3MowhtgUDd/iOM50e9Oi1BoLsd/
8KLcgnSvp8VUcYnQF3VaUKOCnB2L7vvaptJPTlCqbfq81z+HMNUlfzUVKJDD3HNK+5YbeT/A7H9i
bw/WQAh/w7ZAQZGEV7HHm4CbJIOInmRul2eG0s9urIpTawotMJnwnDT00pd5Ps7c7f3lvQ0+XmK7
ce/JBf5dBWnZFdedAoUN3mxcKWjxZhrJ8frGZzzHwAoGQzH/huN6jZ2tAxvBJ7erjWETG6NUQN6O
I7aQly96kgn6Y0Ahv1uQ2fsaFtyoTLXxH+c+oBc5O+Hv8nKx1uPPozIPLm8xjLLNgwJBmSEMpjPN
NtLFBTTnoUmY61L1Y5fDr8k3LYN5qTLnVF40H2kMODfNRFgmTs68dLllxQSbLlQnYsrGwUygiyLZ
M/u7aJ8YcXNr5P1NeSZu9hgrWNRcbeI4jnWrt4AMXgbRysFomiBcbrnp0M7ukPhhcpMYdyW6A+LI
vFSM1bg4C+0KfElnovORzi4VGfnmGvLLTaBNyqCaBJZH3wC9b1/0PqFzs23LkDZTFS8UQD4hICfc
Mlrj44wqOxS5hx9nmIwMaxXdsWgv8PHR2cXdTpQPvHTuNbK/JDFvLdFFCb06WRbWXc3IQziCVUWd
z0j2or4uj0A2tVE2L3FFwWNWh8w6P7Ov5XbOay6XR7lqNckWEi+dTQ5XWhvNlCM7QdpY7e56eIq6
TJhK/iFuKj8NlOZfpoYoTviJ8ASMDiunIldiRpnoNu08+Ci+/wtdMbBVdMU8abnWFlCfW4ns1FrG
j5Ml7NzdM6FTepkKSme80IL2BfoUKPHOtQ9+K8xidojSdbVzZNb+XgIJJGZPhBXmXkwKITB68Hej
C/E3+TUzHlWqql8myZJzZ/Oh6KDBPaneNlQG8NWJb8Ll+mePa51vGU1xwD/NhkLdh/4uisH8GgTk
bUE5b6X2v54lYKziU2gUmGrnBzS9HkjwJxIWHXJ2WUy8kHytBBBbZw8YC1oMHrW3ZBOMsXL7qsc7
s78vE9hqMl6RuShUtVS899NMC6OtvefLTNQNhRpMsqwfFH4bySZmImZLZ/sl9UbsWKna61H3NpT/
pqpZ7vk7saOozZ9B4W0Y7OfzR8SDekylzgGdBGc74N58o1zZ6+j+dXTbsFTu5Wo7IfAyAb8QwjAB
oC3jl+PI74A/VpVzlEHhwrOEzqarhU/1x5V3zGl/Bbk6IljlZqo4vYMrch7K0uv86VsKKnfeyteS
RTy1r83z/slED8TYtVe6+NxZu+e5u5sxMar6NCtswBlFBVTC5mp5jj/RC1F4vdPiiT/PQVf0pfBk
6kahxDCd3R24fpCvrv/FmSRQFXA9yY40HHJ8sL9T8KMSUvoQmklLAxNSdbBcXnQ4IiIppBt6S/TA
sFfmjiq7ThICWCDxeOcto6k0kx4ygJnVrHqrj6ubeamDHUGWppx1oGObIOiZ9A1YUZ8A3jYPowXW
6BL8hZ5dbVs/nDE5kXo8baObG7RSO+ExKdAggmGS4Tb6vxYHjpkV5eDsyn7xYqihNoLW6eHrn6Xk
PZ7BhpYBl3sKWHDkr2XxWknbMc7iqTcg/kkbJN0LzcKTTPH1nulXkKO8XtgRLCI/nheMAA0L0gJz
FwoDDwsXdhvD1Qed33uvjbGHjmQD1IrtPgTdnBisqnOdrktsTVZdgVgY8NTpNToDrdp12yQA3ICe
xWJaTuJFtIrfx9VvTgaCkn0ueAjhxOznNxvub7DkvbLvsMEwDdEL0y3LJyqBletd/dg0nnKTWyQX
LOfIixWTIxzJ0SrfaJt6SamXv104N1C+vhIYXehf0F9FCt6xTs+mE4gkW4jdZNN7xfxhx449NtAf
NLkSWMzLSjLPKcYgktBdwxeCBpleGRyKTv5BguC5x9p7vq5Cwfh+gvgTRUvcEuGtTbt7vyW1Xsd9
za+vQ1LyAyI+AJYsfe8scis7p5bXEpe3O8gqyLcVY/5Ehejrd0Ebk6glTuak7F4MDskIfGiu5h9R
y2DI+fajX2lR2bf2zAIl4zZX2+6kobJodfFbbWaGDeEMvmDWUPq2cQsFBAKefAFqLedZGWwv8hNv
GH1TGKPXvSvJsIBrbF+ODLbrMQCfQlOmvDOdEAKFeK2WQH4TgiDFyOUJzDHMxlN8PHDe/TDVdHVe
s5lB5Vsr2IhJzuVRGmrNM3y5XrvtJ5lWsL7zrozPBj74inmQP0wD1vavJwbjIkPt1WD3XnvWKKzt
UxpVmnvuINlSM6hP/OG0aCoqz79Pd9eaPuLrlzwigi2991hi5W9tO6kVYRVkpOGgBuqBTXOCmpPy
1cJpOjN5sHoqpd/U8kZvCWTJBEzp0BkczCQkMFm2dCH72H6Jp1e1TvwnZjkLaOQfE7E8A4ftcn74
W7pCqLr4jNmXtqEqD/AHx2UKMRrTXW/+R34soH0t2K5oZHkG7mGPinHq5jnT207/xuLbj0XVZ4YU
8rHTpClJ0XIww99KYFlFWzclUx9XqMOTKerG6pSY4Yh/okp/CE/m7j5D2HRP7sKni3frs6SbNOq5
0KtxgIVfY9unuqGHmtmdWZeDla3ezwSgtDkRPW7jzuLOcAY1ImRqH3IC15e3GKa761rRW+T8hGrz
EGFSRF6biJiHibGn0uyidOMvSYqjOw1j1KugjFErBTX2aLI9c7YbwpkkTlErQTIpALM7yqsttKUC
Au0SmXHPOI/5hG5E2UBPM0uwBRLreochmsZMLwJpb6geqHuusDKmD6qlglXEuNDdgtlpkMq1yy4D
VHDe5TajMfDdJ36zjYVaU7yzML0NxhUVl3vSWixizRMIOxpUxQmDhvLE0Hb5mB0Wkhh05Qe+PadB
9CDQVb1ztNSqtGGqpXUykWlJT7W19WtbCw/PHFy26yNnptbCKiarFOlLXikOyVky5UhqJrkScLTo
4Ije+XJffU0oV+f2CD7SlOz/xbW52CBay4Bdbph85vx7ZFa5DeK2uxksd8frg94SFMRJBqg6bXTZ
05yT4DNkCX8QKyw1qgEVP4fGFsXtMTjtbGBJire3EpU+eoc0V4IjY0w+1xLsg031DPR3AHKMWDKy
i81I2w4PNPl68lX3REL6/dfVTg9zGsJD4lhgvNpAbO0hAW3SdBthZ4ZwrhN6l2zg28SOEgqpnlxM
QXIfUqZcyqND2rEsWh5CQDqqcpF6IxJZXv+n3XQtlayqKNmwJe4Ic2woJGiI+A1x/Jeufoxjjos3
qa+P5R0fv2FiZC++rjZC/570oHjKNcOdDK03cX4DrK05RbCyYAmOMsrUbxIEQ21LSPhE2iletjmx
E3j92xM/FJVZ715RdgSsel5jlbCzVpo1Am4/5+Pt4A5QTW79pjUElnOjss9ISML/DztcrBnK+goI
OpeIoVIGQTvt/1elDPpPFPQyEOOGiMvMrrl+ikksP0RiWOQ62olHVR1IVtopoXleGj7s3n8iwQMX
KhOOwOYccgwHwfmx8I0A99NjfVIy5kOSq3AcCZFyHb90+bKzDCY052VuVCn+2jpBa7VhiWCJ2Dff
o2pMY2XmqXYY9+myklWibXo9wBMI6HKkMQK0T2kgVhAqQFurvDwztirN0ov16rmUSeHvBVJWu6hD
XUmNOlMlxJrILs4qiHevW2SJ4gbHpkAFrvKdEejkcjgZJfPpG2CBFnkDdPpWqKmsNRBSR+hF1c3R
K07KyBGF+WkRt7QWQQWry8G7YT2/w/2DQJskQsX4vHcl2yDoS/oCuHPOfMPLVugFNtIukX2qBzSW
mN9Q5PgnHIlz09XY0nXDI6GeF+y63crL41igKJyVB4t1OEOtLAB8DgyuKCpdVMrVF25u7B4lv3Qn
maqf2jwdGGQe5B4h6Wfu28vo1rAPGr7VI6HwxTkwzIGKzGEdauAKyAh6UkWOeUUZzLtlXrCGXrT5
vbEENur7ZyV/RarLL3oBnCc2EJtaPpUfWsO/fcQ8ssZa2BNN5wDSaE1+84tLX3Ui1zrZpH4yI2Bm
W/KtFsV0rcoCfb5SxA4f+t7xQPGz9CbDdAoVgBnDcSGgEh692arAleQi7Phaq0cpU97+IqdM8t9b
Z/YRM6++2Uvo0OwWYLXGJI6ba6pGLS2C8wtHC4xf39Oid6zXVAnJv8kmew/8+eqxHVT3/RFbme9H
c45wCV+8QcdLRsSjxd7XHF2Ur8n9rKwzQ49aTOr+kqDfQIzSsRbcM8CfdJrwWvw2s26OIX6fAqXC
t8ZbBlXTOuIxbGmNAP73vhdbEnGiCk3MdqTwaHOPrBFE2YhRrVPN/BVBZZSmN7QRJTzXrRcnbkH+
tAm4MeBq7UqHJy3sQB3aFvkdXuzC3PeOvE2yzP3LvGYzagaW3V+Mc6q7sYGqegrgYvgH2QqqYEJC
XMHhuSNBcHleyVuaKcUqqb00FJg763bOHJr7sCtLUJ4q3ihs6apirUALlDA6WLkRszNEBRV4f0kP
mMZDmtP/C5rl59/nfwQdgcSOy/5vMSu87MaHCekhtPLFH1dN3EoKQ5TdoZv+0EdlTj0ta91wSPJw
IFlsHeIVBbWmXV3gxYVV9va3CF6XpFe0sVzorxsbVRjueyAFXzVM3DW2JVcWexhqa7SWKYictyjF
vH1V1ZzhNE+iHuUjNeEiwvTJF6FWaJun8rmuMxNofQfWVw0ZVdA+KJj7sJbG77hh45Rf+NQw++PJ
FdCIt6gsPHutZ8htwgmtZ8PbTRzVK881n6wWmnnYTIOyYobqKOwD76YGr6VdPgWXPqNfsVFCu/Pz
RwV54IM/S9HyuKTasnFcVpYYitgFAA2BrmsH4T4ikepdOKAiy9BQLrUj/Fz8QIUaYugG/oFSJZJ1
lHu3Lv1/u/yp9zwVGDqAbezAiOYUQ8qMRCacVib5iPIE/tk4h0L0GxfCMUCDffHx+qc2pb9n9VM2
hniP2EtuDy24geDxlr9GEK/JcMLs3kqrrFRmMWiAIQEBLgMyyXmZVt6aXq7mBIQMddwv2Um8kef+
QnAhaJJwzKmz2X5J56lFHLqOE4daEGgxHdyDukBKS4timhtOs80LVsuEFx9BkolfowwNi7uvrTfP
s4a5lMOLgMpmMoaw1ayvag6IDJXBrSO144vKzXcjpDuv69ecfS591ppkAz8WXcxf5sG3MKHiDjlb
8+R/cWgZyWQQfXWSXZ6UZUT/WZcSt7MFTABmrcJMVqJF06Ronjd2hMxUeQrzpVasIOqkIL6zuFto
7eVcIO0Imbmcue25xiKxBzNApTaPSgR4jPWsR6DqL2TpHALsrytmV8OEFf3nf/yGmYRatEFZTiXc
es/WfsLoC3gchwS3NfAjiWBIZUIUeiPdMxSahNKD/yrjsqufjKyosONDcy58aZKMee/jmubfETSy
lcjXX7tjDOVUfJM7rDSuGcsLVwF65LkDlamG128g8ZTJgy4BkIzCDiHlSdrqd8Xhss60vOpOGxpO
tRK89lS7rrFYywAHfWMe1UuDXMAmy8DuX2VYJeIVLnEkE05MOr+SfgfRUETZL63DGhXM8wGorxxd
bnUEhTqHF8TEb50xkJQ8XR68yOVERS0ZH8H5eRWvP8nOpUit95UVPbA1EAgMCCy0fxkRykp9Tp87
I+PCZSL83o6rJ0UolIqH9omRbQROJsCklZ78jx1MB4aYIij69OIKL5lCHjskdxWC3tqUXT2umxjE
j9QHzNX4nSfoXVSJ+6AF+sdg4fxv8xh8se9vcCKbPqihpRZZdISLLwjbFupZx9VETqic68gbd7TE
7msKEJNs1/PoErhSIJVODF4TrKLvjiOT+WtBG5kOm/Pk6CvTveVYf2ktvNxueA4dKW51p9WaVUXm
uLoSYcIzM91WgPc4djSCDBYx9rFWcXjzreEv886nODfIwR+wLBsYuPFkrqd/R91DndZQUeTBywfS
gZS8tNUJnn+AcMC7rYq8dvyVddG1e6p2x6YLQ9hMAhEKXNpJ4483KzfBWcgcXHkAt2S7Rs9Ho0M7
4Z+fBkEDvWK66kjxZ5lHriuGcR2DuswjJd2XXWvBTx0WIP3BMywaXp9GxNzc+u+dU2Rzeogrzkn9
0zxKxlAITrhubr2oqZ1zpKQtws1Oe4vOpGXePcW4lH/rF8gxINr6qAGA2JRIHFcUQofPrOA06Ggo
kNS4//t4v5qYXh43k/GIyrkkJRCazepfXyT/CJxjAG/cTbXCDkUFIHnslfPFqjuQe6bkV60AsSF8
dJRi4wujs7gyXBfRxOUPXjz0zBMmLwRkKb7Tnoahmo4niWvlFs6QJv1g8T5Mgcq9YZcRxMCMXpyH
Kq+pfha/xPi/XVgzMgFUjojSAaW/RiGYIrv4eO/NaSNCV3M2/ZwQq0t3LGvoMxJIvArOrqMk/SZl
/QEa50QJ7lJB57X5Qqz3PYPbetznfHE6sMxf05UBIoRrK3tg4d98ARH5HnGV+wVRwg9DAaWwOc96
J8PjwCs0rQ1GWE7N8IaDxwUtNxJEJmdi6j/SBUQhCu2OtnhtOJRwD39YOfw/yfDAImpjDtrWfUFX
MO7LFBf85wbYXWm0RZ0inSP0ESqU0k5NBV+xmtCtLJ3N0AQMkRCgrQ807MVwGFhYK2gSfXzuZ0QM
zUO5IVprnsBhaywLk0ofJfsn79h8o+0syFkT2wG/M+9sQjuxDUx7BNDgXIVf+Pjy7yVfV5VGvR2t
PfHO7RK49mzG2jkURy2MVIV0Ndx6VMFoHxywY3ILEbD+JKYRmz7eAOtFb9UFFdvd1ztZ57/w16pv
D4knu4s0aY7RLEY4d18l1UQIwemvjIgJAlfePbn1KV383StlG65Axf3QVtYQmx0Dc5LciamF9Qi9
azuNwlk+AUPYrIUnlt3YJ8g1A2nmPLM2hWPj2yVi6VFRDY17Ez97nunwBT4hj2931Be4nDqGYc5p
JlMNq/26MGXxMhqeFgRpFXlRJyaWvJA4m3Of7deEOyzU9dC5qTLqBMUfF2J9mYpuJ0TuGxiz7Urj
SJVym36Xmj/FxfkloQPoLQsWyVhprfn9pT1lslH1QY432S1O21fgh0Q3MF28MmCqZykQ8rYQAjEY
2RnGOYYIwPZu3yTN57u1h1t4kx63Ip5g6JjqfczSGflfQDXCiF74aEnooExBQtA/neqdDEupxP6e
JVwVrvsNqA0WJEBzhSiKHTQzULYmWNDwI/+A+JbDapfbv3Sax4njKziWouNq5OC09/zCojO4MY3W
jiKxaJ0yRXeY5J/DgDW1nAkdorDpFspBRpO6E7UVIjVh5ksZ7GCIf2vq/AHB60eZYdyn5Bb8jlpo
nW+UVcPBSNQJc8SoPSZGV+lRwYJ0IMly29osfq1RSjzucnhTHN9tZeibjilAcuKXRwH71Lm9sqcC
Hnx30KBaINCCTEbp+Z1WB/jaACkURKcNbwlS8B774jqRyCCV74sij5y0MxHXa4AX1B0fqkVz8043
iDZGM5gRr+qbu1l5RK1rHS8ScJRpu/ZsyXZTYulNtGbIG1vXGSWOS+/T6m9VRCbjeFws4kiY6+QC
FJ9oe+cVqvVs/Y9W+eYJxk3KrB2WcYzkwAW2WIjOy9tiYqm+waiGKOsXWPeQIYeUpzKB4+GSJnR0
laP0gYgo5l0t10Gfc3OAopknITAmcmaP4KjORj133ZkYkuCGD/et+tX2P4VFhK/q4aYJ420Xp1Ww
O1URfT+QCqS3mikwhQW6Vv1+cCo97q894gPD1APYerXmOvU38hUyRw5cVOpwT4FCMY5K//Oi+SB3
VzUNCHaNJjp4kUaJY+ATBlCiyiHNkCLCT17+iKrZWNDL9b+mETEiNTJxZkwvGuEs69fXFs4ztocm
6Spmm6F6wCwHCYSkc4AMVadi9jkuCOQGlT5wbU+Yy/94ODCDq/ACoyDzwI7xIUNKM00BMl49FxHd
m6dF7txq0Of6ZlWyq01s9sagy36h7/kKgKAFuPIOoWxASO4ePdSwIVI6Cu5d7XpM+PqucJyuu+E4
k1ecEFFMI4k7u+T2RHc6Hd5fLLVkW6Tp/0cUQxmYebzPNGNe/wErMTHSqBp+HmWRo5TBrrhYCyB8
LrKCgzqrhcOtWMd15MNhXF4vQgInw/L+S9jLRPzSudEtx25bEzoCXT7KIaZuQO1W7i+M/1rebR2P
FDX5FJsOPSygfAGVurzMiU4ky6GKFZb4S9VzZqlmnjCAPCqkUHyBPkapIakaCb5jhsDG4GfVibvH
sa2yq5caess/zeQNv7qSfqU7ayosp+ejTo32o6tbbBMG5fA5BUG1OrSwd4MjHjvRuCfgAPauCB0N
E51WBKOv2uCdnpADkD7JP3p/9OGKVNUB2DdIaYK+HXaEXeBFmVxzHFuTEMhbO0iR27VprDG77cZH
4rYXGSg5cn3zRl4qv2wbodbRwx9XFoDOchMPYquCBEd61ScHeRr+UzAs5lOBsZ3WOpULA2OHEmty
DlFVloXkqbA8aNzU0JhA9TpthiS/w8YxgbgSa/dz1Vt99Vbt1gmRXvcfy/PQKqJGm8leK/agdRQg
qiLmMT4dd9BSMSCg2m+G3nJrHG1FcU7a4MZf4/TxMMkjlWb2DmoYDCYYnGzhfF8ec2divnpzLo94
SETEf8bSeUlpgxtLotR2YSi7o4fUQiv7ZQJFdgZ5kfY1LPLeGiVGZ1Rem1zgY2PjMF6xvG6z75z8
DxgzfMYxF+OnZBmAdTfkZSPK2U/s9hCzXFLul63TJT89FvAX0GO1npDyFFJ56eYp0A0IdrM1QP4K
+ok6wHvk7+9sgxlhAyHoD5TK+yezVURwr85bx/lKPtLzZ6MxUvKZ/lcY6K3idXn1wUY7Kdka0yn7
EvsILUOMSKpq34ojnWQIIAm4F/qveoGR2Q1GjaqeqfdvJTIKMqYYAmsvkpmx8n0+cjPyJ7od/vOn
5uppskrRgQ9eB2US0FQ/g79REKYImmnV+El7mYG8JPkpKbhxpybylOVxX2fjvOfn/fWceNoQtB1C
fBmtTaC0z6pHsO2KlZpLi09EJPuyUBe48gi/86gNNkVOiq9jFqqdhel4qygke6N+Ttj9jGV47ORi
w8n/cfwvX9Kt+aRSux99nm9DSuvv8rsrE9RgCRq6nQqYXGLYwYuqhalp7R63VDIeEEIUqsWPgnLy
5IHCyIQaTULFYQZ334V1m6I2qWggSWUwGh5OanFkPDaRgm+V60B+MYcAK2gZR/5bJs8EKno9v64d
pNtQK2/JuXvZupaqASylYq1nmS3LVGCgLYPRt6+RKfYhE/SUWpGs58c9D8qrWETox9YniJau/0Bl
SjUHX0bLl5qYzzuWKdS5SAO/BrELJu6o/WXjB6Ldpr1PoS+JGd0t/EuG/a/WvEi0DDgwUtotG8/x
bZI8Z5OLPC0XizRAHX9Sc7F/Ts55R4ryfvNKQS6cgVUxvzJFZwfpLAhpoLgBATQTlqPqAI7LZirG
PgPjQVlBx5ZZE44mcWS5ANIIRFItUNzowjhsHVXNcDGt7d8E6yJiCFacoWMe6db2lwNkgTRsvznF
lT72oSScOvoCaVQiQ93Tw4BGtPEU8JNQckjhxgER+9lTqW9w/tqSxDkZvImHklJ+wOyvbMutk2T/
815sX8iZjZwPVyklSKkPoHDxFtn3g0gsNOE+n+6ZkYrDQfHA3faon6qgwFPgIWLbj0w6Vwm0oWzm
QPD7vlZDxSZ5OSJHVy5dXKn4psraB91UNhe4wcb2co8fbdCijSZgDn2VahfLYWQI/+KJSJVOe8Vv
2cwdultE0rUDrOuvvvuU+XygabDk8vhbsFuSEoY4mfn+h59aYP0kK8ibTS8vny/X4z/EA5kqKFJx
YSB6HO1yb6tJFZALb7ioLDKiXXRpm7w+qddiHQcQmaanDrUzOcGbKd5xqraEKN85IoXX9LibEfnf
U2tSLwqtgYs4Cg5dDqx1YUQ2ptNQoYJzUImyBZCEv5y+nE9uBxbOMQA02f4ST60TajyXzo33DYie
7M1DoKfUDgvUsNzY1CRjL6P+5UPkekZ59Zx4zBhFEuhanTxldbIwsVninr0TRInd5kNeSNC34iAH
bF4A41CZGq9yxB1cAhdCPn9+aOZd9vLCez9t1PtadBG0jOaB7ZT0lx0702jP6rtbnWVfn9a26pxq
XxCUGMX4+UAZ+v5xeB/aKJao7/fEJEqjvgE81UBSvGtZGc8tHAhDabJuYNqj11F0g+13c8ir/kGu
NRvvlFRCZoMcaWW6mwwVZciQPRBE2oJmUgpycr2tVhi0xK5irF0VukcRbj0qHM/5SiTeL8bDHkm9
0R7J4YWMn5Fx7HgPb2FrsLM+c1Ah12B4DxmiXPIs+0D1RXbXX8Z20EJ/85ZVoV7hm1r3Tqyt3kIm
uVz61JXnb7hkZJQ8AfucvS1sWy02VASESVblDvVpyLmDShGgKbkQ5NaD5iZko9omUlxKxO3rUOg3
/HgMEs/3zHpuio/4J7OlW7U8btMwOsZAzn0v32wXAc2LO8NW+st6E8ZFocazll1CWyO2eRpchVlq
evLbT41gcSG/cIx5b1X0WQERH4Ept/xbrOwBhHZSshtMy9yXpZP6bXqV8aElBClRnxfsnylHyUSI
GQ3K388iJPs0xmae3fpYPV5/DWlm4PUSnj3F8WfrTNaoMtoa1gnfFkz6fpxraPoxQhtyRKe8cYOQ
PBDI/8uw9LIzlj9l3mLREKTbBr6LABXTv8f61y1AXd3EkfAbeO184O0VSiWY4tIE/2dhaTzYWddo
3nCDvYhI7WVFSWAdNV72oq5YW05obHujHo/JoieLCMHEfJBuPOUa1L0qsZOjxviwxwTrNUb3Nyo9
BpT5151fwrTCHnIEF69nO6sseZglr0hflakT9Mwdlr7VDWeblYZuyRWkA64Gek2Tk2k3i+79vV2N
mrCGdvjs3azTQBQGOc0BH9WcgXYQknjVMUs0wMu1Fz2XaeGGbZjHFliaxwMsyZGRpM+3RGSLjHO1
+DP3d9LrGiyAv5NZCkRPBxBzAzYb3fwbpt9+bvBjNkgDeMusaiY8ud1LfZyxLPOBJHXVIXQDA9ne
FR6kSB1Zx/+ppTcrhaUMwztU1h96WL8nEEpxA/zXC0m/SuNbqlHsMzMFzmPuEI0OrYLcOjKGaB0B
kQqtwkH4qmrsrgizlHVQZfL08Lx7NDzmd0mjgpCu1XwbVhB9ZCU0AGE9emzKUVxAyXEoq2HNaxaE
+8Ce0L0oPiCd+WiCbwCHE6sw5UZDTn5JEUDxYcq1FXQXftiiAtDiQSLnsfRQWuf+4n8DuMbXZtN9
Cy4WHc1CdCwLDy6A5AYR/UMww2prz7vuYLAmli/AhpAp1cIIpaCiNi0QHeE4MUaffjJkYsPm/+5J
OcYaxzkwuXx7ysQMme4IT9pNqj62Ts6GiULm8eZmKRjUjwTNdKdhhMtKku/zOXCWmCl2clUMTwtm
FXBliUtENi+qIRQ6bHtoizhBuoqMKZQONjg2fP/A17SNQu6w67U7uD1GoTdS3yu9ubMZQisAe/xI
+iQXxWjNtJpQMFNoY+9kh7WAYBfsM5rkI+y373TMY8ANk0uckWG3NncVBnrF6ke5DbIVdMlN4HBW
leVeusbaAHaSEDbEu7rSUs1Prvq5YJq7sfRWWLpWcObYY5cEP61py1j/2xksnqkRBOPNxtUJ5Yb/
KQ1oovNn0AGJcAe4o5BaRaeJKBK594fdx2PPmkhv5wI/h0ldnW6wwR214VI2vS9qLmrQgtJeItag
COo6XYrBbIsl/RA38c4WVUO94qfb/N2T+zeo9qpSUQoqixWJM84cTVhMRrkskGbQtK/9x6JkFR7k
Pev5t7hUhCa7hfIGua6o7H7FFA9vu/D52k1jtgLmpHXyWhM+jh9MHm3880kx4F3R+wXtRGL4HYj5
wNuRgCt7to4IvIkjc0SWGD+vjYT3eWIMyvV6H3iLRe3eJJGQj0U5qinFGfw8fg3Xhe54t5J8N/ah
R+8QXsJXxSEzr3TbT8QLbE9e/6rp4JMjkG4UFHuY6fb3Plwr7mwda68MOwCxYAkpsYbEa+ohEl3u
gL1IjI80LuAff30P3PkndqYqIeiAYhA5cHUeJNeokvsgA3l+PQYKWne3aprDYJchZkBw80jLz2S6
ZIOXa1ETgBj7sJwH2kHs/qfcTT4N/sP3mxNiNf6emUrtsCNiks6SeZpfauymd6Ys2ODspkEJF4tz
T4KoBIxYC4EtA0lLS1687oIO8cj5gIyNB69kyY70eIB85HO5ZfRSFy9LNgDad3C05pWoROBPOVdm
noT3TJrcHd6GWLGE+zkQVnD0VgeuSfNhBd5vMsyv5AmNukvIrQtJz5YNG+ZiODDm8oUu5N9m7gTs
RqJM+E0XrRE/nHZmq1f3lcmYPFH+LquUTwbeFcRXAC12DUx7fc7YfEvQJnZNj88LucLdoKv5ur0X
fbp1oiKvfnn6fn8eErxIO7xmBrU4u0OHQd2l72uY/UDN+Bz9MSgX+BqoymCpKdvFOwD4/1l4UpLE
mqHl+beCQJqg3Tym+l4q9hvYQ77vE6tAxVMrWHBqjtu/z0HS3ftsGR+zacmExudrFHnnTt0dQ3/D
/kGAVkWpm6t5UtO9WWpf+6SAHcJHmhmjCGsJIr5P2vfJVM/+xIri61ehEP//vvW/mjq2BT7gZLYq
PXWQT05ny3948AOnTP2yHCmqKP9boiSDfpr7P/OP9R1ISqQaz3BKrXuJfpVtdnO7/1D8c+yI3nKn
iwlNJFEXe5D9rDcS7e61ldMRmRZw6So6DF0LpC8d5x1m8hwdqBP/aBqC7lNFWGtGbaqVCwcRTIAm
JIoGUYcnZeMYuIqvAXuqAVmQmnYdj80J440kYTRLiBTT01x5CAMnrGf44hqy4c4I8R5yGl9rVl0t
zBpSr3hhrY61ddsQ3Iv+psMAYDT+J1RvicFR+hXU0KssXmVFQFimB8ZIvKyKh38EyumJDtquk/Ct
sSAJK3dyeviL7Z2nL33mBt59FniVJdBC9SCAzrnEpLoqWuJS53Jde0BMnMaQhaYy3qCpS8/E1Bxy
X7yOhX7tFYTpQXtvCaFx2OnYQNzLJNN8AirbF6KNMOZoacBw8FrJJDYGWi07wyMfg38m1npPBE5w
wyCMIKHxy1EaHuhDvSeit+QmKdGeSa7Mhe4FTVus+Oix/iaVqyNqWrQMkAQkd/xMUzwcmnYi14IK
OEFAPR8nIirdosVUs+LroV0C3EgQw0ynUx3gnI4wrqEdmBNeEkLuD6pi3zw4VN67ogEWuhcCmu/4
ZFev75KrBhxmk6Qe1U0hfXmn1EuQNOoYUJL4KyQ8Cxx5gheWZ3/Qn9ezvDclomqimFDt++p5Pz7l
pAaMB+k7mOwhO85uYCn7SsOxYXVSbIwpR2EFWo/D7MJzeJePsxm0ZiFyVd7W/5CqYZjKQ14iRkal
JI1QFdULyDsmixEMGYcK6tldfoCzBFIhp+wQw1Ev2TBgz5RyoeHwIfJywPXEJf+cbbMKFLE+GGna
7zI18AAd8ztA16tzNbFvYvMA5SyT/JB2jaVl/sHNzL1E6qPcmUFBy3L8YuSuSGYKICi/yNrrpVmS
HVJfgydfXk2eGd+JhfpzDQZCII1tO2+KHkRqZKBB95bNBSy5MaGL/8hjgr6aQwlhkXscvZIttaQM
9EP7wfmHjX9gWK9bQrqGvaDfgIdT1FAhTexDTuuywFXdm9jxKe4xMKc5Lm6cxDZRAk6AXwmZV+eQ
ojzp1xaS+W3R7cUP7HkPdIsozIqQ06uvd/fQi9w+RxPKmyQxCmXWzKg83WvfsLh+ANAj58uKtq8u
WtCReNic5ldSIXZT6cvdSGEWR2Vjc6w4J9U7uO0/I8w/2KhhT3HDXRB8sdB+j57AaN8/QYA0lgwS
nstXVF2QUZo5D8slNBByTX4ZZ+Q/WWW1tMBU0og54DcqjY6ofxYrgczrJJVm4v7LFZwvTez7VVSb
lWyd/WKLxsDCIrN50rdX7Q8nX04RK/0vSjCP11ic1tYp+olV1oL8pjDddhSNf+SEr9ua9k2QuSVF
YoZQIlsY1HP5Ffj9ZGTcGKnO6GnhNdCfSgjZ42o4nfajwqqr61aRUgAyOJu6wdD3S1kW2LxGJShe
R7W5Z+xslKkW/sYxZGMfKXHQ4j07m6PYktONxHJQTM346C9kU6LYkVMfWb07WmGsca2iFqVFmWEX
COcKlQ9Xfnp/qm9XpY8AcD2PUhrTpcUHari2YrJmDt5/hgp9BB5u4htOPYHr6qYZJnLjZKjbl+dx
XvjEIgt9SodiMRaSirMtDo9R/IaBkDHjTJVS+MaUHp23cX01gpQEPMLus9EkKnB/WXlJTIX6uHsA
r7htftpFz/iAfTSNZZ6KZhPBzXme5VU6zsDZ0MFUQ4Zq1XiUfDdxSuyBrvRMbimVgLAmYi1mAjch
oXlqsHEjdMsiZNw0jMGvUGm9VET5LgDBivZ6is8OmcH1BALBb+mp7mMgle8II9KeHbnyfDQnJc5r
RJ+2ATa6JnK4cWhOSaMxTq4NYNMTTsiU41jYp6TUjUFgsBfyjJowQJIEEbSXDK0bKHbjYlts3c+B
sZ2wRMz9aAnJzYWQATYIs0Gom3RMSa+bP52xW3/dIA0K2ZeN5TgtzF2sKizho47hYntpOZ9HT83V
s//KSYaXrYLbY2uDCu+KCqgICZV5buYwxQ6LeQ2ENBaMBS2RstMA7RhhGaTYqrlWdK52DxeqkLSr
MaZcsNFMM2oI/+p3A2JkKOtNH4U1kpp6j5FBX5yG/3XK6WSPGXwBpRR2ScVsma0Y9unMs3UMutmJ
ixgsgIZUAqYV0NO2RQkKb+08oBqv1faruPYI5opAHT63MaF2N+EHRaltlq7OlOltTg+1KnfOKDJg
zLZ9vSMPK53wItueksu/L12ZiSbDTDumyAa2kE9z7HiuPGk4258ERdCJMNnrpV7N+ugaz8fSUqsO
6pbFCeBrx5rVfIeqXp8RhJL7hvKKZjltW28qmQHPvMmRNK0bsffiC8vgr9lSW4uSRr5Gk08IhW1s
26c63ZhuLRb8sHF2xA/d9Z8HNpDIgbUs4awXLyyg3BAEB9KgkjQkUFi5fgrbHVqSlGqE4Zx/UNzt
YUnubW40wACImIncebWywk1EiErpSN7dy4mxlOGffJpHMEucBP8TN2SOOzyAT6ziW1Zew6BNZ0PH
VbJl81O8s2G9OMe7fpSUFvkHjQA4xNsN9B8sZJHSTm+9RY8putaUhDwKVvQZnQvD0+awKoKvZ+t6
5by0HaxLn93NSfhgS6zMTqpP7g7i1pUWce75d843xTnw/ge0opMAPC5mjWBVquCUQl4gr9SHsSc6
XJNXUrhpnPw9khOg+AANCbIOE5UoTueWH+BW2z+Loajc9DbvrgL4p/OZpby6EW33t2S4LF8HRWVD
pOguDjXyO+DEmtjDxB82qOSPVOSbRedDwXmfNxn8Y1M+u4K5XpahB0BWfoQfE3PTM2OAeueMni7E
d9gPkUTPEb32u/vEvIyD7sipE9NtIDxCFuL1XEpNPw6uKvv80oRqQoTvx6i0rbbntrc5CU/OqyQn
UVYvDV0kHm8PKdO7bvNSQ52GkL/IG+DMK0MXZYX4EgC3hf7DwVEMv+lsgCujNO+Bc6CugSorxW42
2HKhv8p2QXLbDISsOkC91r43kXT/wiIWwadF7cxTk99CnAYCCsvJx/HdEjADPjltk5D5JZYE3pPJ
OwQJZVSU3OlRXG0mB54IZ73YdZFKBAtUsoWz3GEgoBW192NVqLNeeOs5WiZNony31huPnEJOCwB8
ZXyD2Bkw3LJqWQUtokTer/g/bSlQ9x1Kcuevcm9zqyl33iFEytMW9cmu4JK1o+XPehcXjKvin5q3
l+7fJ6yVN/Y4Fz9aHisRyo1fWGIirNhqAnLvTBc+3rC4CnopIdUz2H0im/DTwWuCRRI/pHaDzWAr
Y+UvoPc9W3kMwRneSe8ZYhIa4Rn0nuDKRgEJYAEaQa8Tt/MbQ+u5sk3S1kUiv48tZo6dAT9fgD0E
sH0E5LCyDSKQA+YtNmqOe+mgk29gZVf9Gtu8yCj2iQeEofEpaQHv8SSwRux/XqVWBil57MFvFWCk
1XWPRoBo3YqQfm+PXRXZnSWg9L006HzNgoTOSsGj2VNoZ+pdb8df+Yv3EWGpjaCaj9PLhGf+h8TN
31zCxRxqtwPLlisLA1Q7dTw9Kwb8cKFEWMK5c2dVT2F08TlzBxmRvCoibUpPw+50/IxAyh77QNPR
xwrdmsD9x0BUmqx/etj1FXN4yLCuHSPwFiSCVt2YxJ0B6QFwnQhJnYkXw9sFxuwMVcEzU2j0ghRQ
ch+HomL3hoHtkzvicgjUKEjH35R18BHCE9wYjvAI9UHfaB2KyqioLpgKtE65soLfRYoCq8ETiSNs
85Ill1z7B8loKwu5TYD4ILyNjRgn60RTEpFhAJhWMF4P9dYSDQPYRtC/LPKEdrWRt91sXByxAkQp
59T4WQIId9F09NVl+dmi4Cv9db4Mgu82uA6abtGt2vN8SgNJ49z/vwk8rxZFh2SxIRN0A4xZglaL
s6+rJtkx6g90tCogY6jm+n7tmKk5XVTYmih91YX66wwWtEkHk6fHiNlGA/r6JqbjRHrxhIEVyOLQ
PU0enBUnUbGxy2R+PB9TAJvLxXrXF1kZQwwLBycTgtxWhBsPsJj67ug0j3RN+nmg6sHcFWO+/hl8
dIEn6YJPnwxdS4KpW70v2aw4EUEcEr2XKGiKtcK8kYAPJraw0JNERM+/Oa9ewnzqoZqbcVmsmKhN
zVNIb4YWWkxTySFlIcnj5oGbcgPzR4byMGGvuh4/x7AqNIx4cgfyY1Pci/GWX+aPVwfW0TPo4yA5
XgjH68jcdv9JbfpvadnWZrxDD9RA2m1F5tvMjbRWYEzeil+zPJFFOdpAN40h+tcAy48KiyBdUoiB
a4YA57DEwBK/uMK41k18aZzTtdBSXP/de7ihb9xr3jtma+W6oQii+Q4wc4oFYOY0dIJfnlC82MLP
9NwV2DPUPE3x2JOPHclTKRrb9B+jNgeFlCJYywA0+JNEnB8wYQZPW0mbrSw/yMoUkTO5RS99QZ9M
jDqVik3R9rbzO2d06FlSX5dBNY2j3hoD8PGynbESso1xh9Gl3ysd5c2YXu7YEctzjI3X+x9AZNYq
7xBFwL7m3Q/PgpJAHsGMoWIVLiUoPyzVOU2tbRaRt7urjYJWxC+++OIuZ/SLv2KN8IufPIt1dFr9
4l2N1nb2Vr8hg4bgKJpNYGcu5BFk2bU4Yv9+6Lo+fX7O3vOoy7xD7jgmw5BMlxao8m80s6EM7gdj
9gJbgvDttLQtlL8hGIvgeRGssPzTnsI7BZ1UXdX3+fyuEPgoiOpLQox54+Iwq+xGb/GjvSkjlOjy
iGiBqqg6Z+oDBVydJTPw4CnKZYyz8api9JljpRW5GRbMD6WmKX3zlkowJolL/4FwlgPNDxkbLPCv
H+uPOhspNFgrnEGS4hxxTt9XZ7Ql9ZKIo8oaAVlRx924aJj8SEKuCxS9ICGIU89qgBTJeHi7yInI
Bhmf8t2lTabTnrpVygmf/2hgxvasxeXyPqrC/IuEio/y/ZiJi9ssmpEbwe4XvrQOzFL0E4DvdrrU
s26OJkVUQ7fgx+fvmyl7rEaux/zUsOLBLrVa1OI4asrk80Gi+aJKPXMKHn1d0UaViPC/8GrzJiGV
MBkvuoWQu3Kj8CoEMyY5VGfPMn3DCtgg9CWtEHUpThcPRBDNaDxB/si5T0UId5YBvOWuWnIc2vAY
+/omnFY0HZALj3QkrV755WUTsTDcDxgudOSd2K+10X7ZQEqE43lQew5P1g7Hd3P4A/iCqNHEnfA3
0FRPp++LE3C8AvNw+UdlkuRmSbKMgHQlpeownujnThMDVTlw4/PQWgGVpUSCP9RDHIx2ztcrxFl0
b+s4u2l5pRlGwVjIHg+cWEKBMkLqXAfVQCCnx5FmIn84pdtt+K/ada+2m/1hiovd9Ti0Anhz9zZR
VMEDuA8D2G6nOixZ6bYx9Nl8dHDnmoCEFbicPdJQ6k3Vzz0sSm9DZ+wYF1YZMC3amV5xjlSU9A/K
HaVxggwwdHV7hPIt0MWtKJis1u0rTyftpdrHrQAFwuyt+H4jI7Px0fI6sS+0gnjrG6tQnbezGfMb
HO0B0L6sJZNmBGC8kuT/xBN864aWOI020tdNWc0mN9y1xLGqMYW5l8GKfFv0OFnUT1IZSZeJdJ2c
4SfW2AW8PFdgzLomw79AHn5cOsk3m0dbQPBs+Bv3CVQ5ugp1zQRzWMB/0DL2JEKPUi143BSLPPY6
Wl6zkuWG0ZNdup8B2xBNkkz3S5In4frpIJYN0VP5D18oLlFkXGuHFqiS0JEOzHBG9nishyetGBwc
Yq65ejYMd3W6y1S9Dg49NqvmNl1gmo4bAQjiXZjMqpYQVkPAhmkK0M1CYamLwJafLftcBZ6h4Dnh
JzZRMn8aJ5dijHEAsSar5kqZBZ7U6tj8RCsTd4HtukylMj0W5cdQ+uZUa6+DbafAfSOcqIi8alnT
EUMN+lL8goFO9FeseL8AsBmJqHhTptSa6vFOL9bRrZ3qtCuSTbBOHdHR/RXuOFU8BI3cduLRBcDW
H+RBpkHI3kuCl3B0MXhq5+wrCma3dg4HH286zm0fF80gC0xuiAtGV7wJMKWOHSFXmj0T2uh9CdTE
eiIBe05ucxWAaVsJi+L8zznDSVSwUIrLbPUxyivFFr3aVkpTx8PiaLI2Zdw6NVOg12bXGgcraM6n
/RpAZ0JqgZb8ZDQ+T27o1fx6gO674EY/6CMVx4rSs9L7KhKcSRb/XfkWuuUczAqenaIp1ZtIPiWy
KL/Dd+bmian+yLuwYQQWORx8VetDC/aO1o/wmN0po6it+snx/chvZCbYnmSqzmFnWgerTVrebV9T
4xIY5O6LtZ6kF2i8+88idk30oi/u1BFpkaHaN/VJTVpoKlNPEIs7E6hNpQ3OgigUQ8i8fSFglvae
1CE96Kz1yTFMCJbDYW1whCEO6RcM+4YPmITKCoNsBlbUy6Msete09zLHDmwnMMdBdztLLlPXEGdr
pM2b78kxK8QD8wkgvnwjHVLqn2JSenyKHm6LvqiH9GZZogrnfj9f4OdGDYMPn7umB5j7Od56dhV1
XFZrsI1PxoSZzfMeesnGholNHLWq9qSez2D2mz9QTTvzEFia6aE50ViPnvGiJdcuh3sAmhRHrwrE
tcYyna1fBAsJuz9mc95or28mQTSt3d6elFa1aAp5GdZMH1a8oxS2UmY9885q1MmHPeCJgO+s3NWf
bA1yEpBLgoaUBe2GmQMf89XztVflqXSM+sFm686mFiABDdwfebg9UEg+NW1RaxbRgK7xIsKyFQZJ
7QX02j2iyldx0GJTA7999n5STF1HzJ3ds/4R914d3NDmtPiDiEwgGhmCjbOtB873mRdHtoJ/+IwG
8KWa+m2k0GvwwFkpDf2DvgQr1hyjWYhlBbEuZzL3NSD3baDVIWZAsQUV2kDSBr8EHENqcb2YnVI7
0PBEOdELjU91W+8c3GSnrrXyIkgzKBiJG5LrqpareyW5moOB2NQMyWySwvsJy17ss6CP2pdhiPVI
XL8i8XBayPPtVM3ugGsc9t6HZb4+3Dy2QaHbjj/Yks+3dRLhj45JKSIYwdDjQ1te+wmDS+TpXgKF
YhKTPUe94pYlvWyVvAE680ot+qRHOEdCWhTT/FfKMka/uQfGuZGiF/Cv9RGZfeJIz4oKdPfg6W1z
iC2iptnl3gIvUQQc1ZQhXFEbzG5MUqKwUuBkWHIj9dYOn8BSyOc8gzapW2Rk0YyWJVHP0NEDvOnC
UT5MF0S1qwrZSHgswIabKMKxjlAfIgPJ6VRaxg/jSgeavA7RFcyAOdbYK7hMb3E9UfbMdUJLQxcE
Fn8qBXNodmai2DXbLqzt1G5+So2khI4sSxvwkKws0Cea6e6vcXcOrYnCdZH9vQedZwCTm6pCKRdm
v6aEYXWzMy53hfE/qcgzipsefIllxiWTp0CZvM4hA6V9QRmVxjyjGspkBBqWB8OFn4ssecvRNzCs
FyABp/zdHkoERSUXfgwD7DBCxHTN8RjF5mfSvbvaYErELzWofVlpk5UBrNeR6oOI17u2N/ZiSR0R
GZ/VCQneYNpmOlXGCNZJJpgQtk44rxF4RNAl1t5wghSVQGAPSGR1e4xwEBB5SPtOyoJGJ4qlDyM9
1P4TiaYOgxGNJHh4R7GEABCmFY0fVuqhJfGe9PBo5IRIPg9lpLhgOSzgOl2K36RyiNl3LOjrXsKb
kRMeBxLoWeJq2Gr17z/J0beU1ov7GF0k19qlc/1utpohM4aRo7c6JeMvEhse8AptzOqugOm6yZeQ
hT+jbE4dX05tIpTY5AwUg93/f1CbWR/WMSrB+uCTzWKidujffSlWiUt0xGYLtTcipl0U3JVhDyDq
ZiUzWOPgMI4ClECVc8RMa1rLG+cQcrtcOY+Ev3Pt2qKOKko+uzOnpSDYA6l50b9gijEUvjGMJ+kX
CxZn0OAF7n8f54gbLzrQNH8nK5UyFvlqEF89EJrwqYumjO3y6qSwp/B1BMZQZ78/3oS2dABr5hxA
PlhxUDzEGSCIqQYYkJ2HY7r6RJ+7aFuMZ9YEVQOfs288oO0QS2FAmoyd3PKZhUfkDw11inj+ZYtz
e8iRCeEIu+CbR3jPElerlNpBf3pWgWvsBcEyXVeJgEKatIuay2zZAS6MFFI5SNCEBgA1SkSXdvNV
qbXYD21UfLsrfgnMlng00N3JPlW/ysIMQx57tQq4wVp/sY3bnzwwlE1sX//4syncWf8CT3Y+oKxO
AUoJZY5K3+0RYvWTtLxJwvLp6GKZCQIhito59j7JdEY/1lw5zgSzj3Etg1zZYoSGbFIdvIbMqIGh
oa1HCy8J6OYSDCLq427G2tZ+jQ+KWkww16G4TRzjXlGDDu3X+9P+/rTQ6082JcUi8RKztF7etW48
oYb3upyDZEsUWsNRHP+qEB8EZCmhW86qtCY6LG/WTBydCa19O/5iZq+/Ac/D0lSmguB60Ndmwvmf
TRwTulWHMTUd6czLD+ciMO8QHeW0ll6ED9PpUxN3WRGYgrDy+j7Dw5gmQCAjl0LvbdIqTS7uO4DT
eLFlDWaMF2h4koaSR/DsWSQf0BYRSzYjochnIYBzS9emWg7dzLcmLbZvxEPkOZuVKLGFN+k5qyFw
L0cYyVakn1KXiEaNSAHW8CiTuEF5iqzTrht3JMTKvD1uxOTS14Ik4c5BtxJL+MEG79SuFPTbqp00
70zYeEjmOFFdIVoBmbwCRVimbNcxZeufBlQFsCfDoPT0MysSsBZSmYOqu3zj917J0PSiNreAFlnR
BclI5dFj/Dv4Pvj9Jjn7eM2law9RmG/jpFPk71gw+9nOeECz5BwSpOoXN26uotnkTZmylUR5seuf
8RME8+7pMmcNRGS7SNuinjb5swbdaNohHlf2MlrLCOzOlv3pcXGTpczyXcmEvnWVJ+8vObGKv06v
Jrd3iLLkHmNjYNO3AU5i+nyD5CyfKR3yMUkM3+rmIBA7S5LRm6Ad0cJRB8EBC6S75uecNf1oadz6
9c+r4WFn9VeAu5VLSL8kDXbo8HJzvJNcYmABJ82YafgnBNnaP72EEmJtyUhxUrKF4O4k8OAwdXjI
iuQTGAjb5S5X15ecYNKaSAsaS4EVIo3il4uBWRNIEYOiiJb6R20rQQ9EytM2IPgVq8Rpj4eSiJOP
RwoWgVEs+TyGPRrUeUKFYNuU8qT7x5vywGXwbkdXg+z+dC5MzlKh2A5y98sTQG+UEZkIW49ttVUM
jMiTUOM6+RBVIAbSu3XbHis0g6MqV0nN/9pIGdPrXIx4UyCgulwWs+sKhyJbGi7wOoukchU4dLdw
RO7yWY3suT1qkFTzd/4wZpCx1m/b0orx08Ta5gyIhrY7xmucgJBLiUTNXkmIztKBJcXjZpHhc+rS
tf70cofmFotH/Fip3Rp1+yYMx/d3k8LLbbv2SeANrkq3su+uHxvEQ3cxiQhavr3+ftskxiLgq1ET
C8Fj3jx27cNovZNeeJpmpbmXZSW8yRq1mNkgV71lxVc0VYkyFXCatniFzPTa+pbwlbLrzNZJihyT
6ji3eKnx82amXXRyhNFbSCdAy+1LZ5nThDpmrxnxlVB1/tTrNqFLJ+sAR9FAHEfS1Xq9PgjqdNy8
32jLYIX5ll+WiIexZgAEOUaGg6HHGxNrbQyNXSjhA7hDWrVPaZ6ZTm3DgnV2SZGRAP7kq6TmgWdF
tBZKFWHGCbfsqVI7wyW73UHTpPzoSrCO/dN/8RXfpCyAvINyTngzRSRXhSsoCxTygDdg6+LZG0JX
8yvOjfnz047zGIs59Fybpj5eJAMj22q4+EWHaILtdq2H4JsFHMukMmeasglrLZL/TH/n2EvebTNN
25PoHHC0jH3rO6+4cwzYYKNXzioQO3dMCYLjb9njRtDmxnkJ7u9NEP8wMl/mWwMa5Z2W42LkCx08
8S/xBQPX20xG4dYaprTxmwkgHeuz7hm0JbzFAc7AjEFq7q4/aCmsljh8okxMgQKuM6tdgtaNxR8z
/8qmMVoYsPUYRUrfFb0AljWOjcF6WxWPcO/eigtSKO8nnihsT8cSnMyyEGilosJAnLFrEObp/KME
XKDDvXh39zd5om8dQKD/avS20lYokL0AKCAnaivoRGBUYekyvgpaStdMBdxbYKYuimdEENcwQno4
dHa3sA5pS1mKkSnecepz+tzFhk4XkaYwk1KXQ6FTcAxPCWBdMnA8e5zBxAzVzT5jVnUlS2RvA8hL
bSXX7fWfcWDaJH1m+CSmo9gxdPTYstQ/GGMhBO490qCrOvkKpFnCLDPtpQ6O+ORmR7cgZjm3fzPI
ZriZqykgOQrsjUnV77fKKuv2el+yy/0myH3znTIFDvFm8JIKLrj0qVtEYrlLAwGSo0cERrtuD4Rg
I3cwpUVy5I4YvzefQhe+ANlsLkOYn5UCPRQJMfAwalv4AcDfdSMYFPvF+YNK9VhIuE0CeuZ5xVuN
QRt4IPEhwH+dEbExl8WzcqS2G7g5eUARnxIXJYGpzZp7iF4Uk+I+FYbQCAjzAOKyMC66DzcqVSf2
hMlJlhbcxSmdbHSe2d0sEOakXzHsuHH0YPo91A42bQMTqWMTaHUs0YikWrf0BksYqn5kU36MSuKI
f7NBx6C7GRkzeSG38fk2eknrZWsgqNndX2sKufAsl+XTNnxr2KcDchwmNn2ufF5NaI6jlBebZqlL
BFP6mKCG+83I4ximKbWiV7KPyg2VU4HIFBP0FWrlW2eGmdHTiXxv+liAlWZipR8eAQIQnacdkclw
yzwE1lgffaUdJ/VH3CRezVOUSibkrEsoITTrLDljdcjjOt/DdsYsTCNaCCSIN0+WBnyj5UQ9MCMG
V6VPygQGJoWAY3lHyYxDjls2KrCPIRKgQfI83rpSNdD50+e+QPcmawdyiWSGqqTmFbR/Dpfkhglg
dPOnxQnRE4prLC+RNfn87PGiHlWfGAyLE9Ybm4Zd51FuFd9QuJeN9IKr+C21ZtyxbgheqKVl8aIB
fY7TZEiIHbRATe1KyfuaHj+N5Dg1ymlabSCb1lEqbXhsMXeXA7DPUvtaQ77pnujtZ1q0knFj2580
t6mo2SSXAWtjBX+NWzZUICMNKz+HBNtQNQefSkJTswTadVw+FYjoUeRIakLP3BP/28r3eViPHhci
Q2lPL5zDSC4AcFEAzpHBRYKzmLXwKYaIGYgVuZoaNumZIaymx6H9PXHEQW6ekYp0y1nkj8UTKYJ0
IBlazCUuqBbEKfLCfvgb5Xfx7c2OkC/BEqD18jvnO2DAx2AZ/nYY5BITtzkkVuWt5wcFwpkS9dVF
6/rYOtZpqSqKvr2ye33NaShq/qTvdK/wWSdx8z4x/WwFwHFEMtY2e86swYkIxcezPYRcWQ1Iggxl
n2ZDY6ubjeNzcmN76I0C9Mnnw1MbX+cSXeGppTc5K1v7/WRH9ecbb8dgMys/r6QQbMGNKOx8nXvd
YWFKek7dQVOWsUbFkS6rIGzsp+b6b4stACk89AtQ6bjuE9Jk0v4/7OpM1/llXvHbNMaOpdwoRm2H
AJ68ETUDWmTOS95d9Htgn/yBI+rLc/Q7dJQLMP46Ph2OSN2iWpIeKUPjlnRqCAZtG4gucT8tqo+1
8rSScAgDbKuX53DaAnOHPoNX/js/wwvro67AULaoQ5Bv9N2dCg6qjYb3Uj/QTuCjYGexx8Ds0pw1
R9kRSfzUzkYU4/NlBeXWphYUIks/yM4v7NDQP6btLmVOIToeoHgLjRzOF4PWqJ1cD3ysbL44AIm1
2iHEJSlR2G2/BpLZrSFtY/C0+hdZ1duuIAI3pAjjGoOUqmbyFCTf0NY6odqMaEpp9x1qZctXIWmK
KSQwGLxBGG+m6s1U/jrfE8GSVxb5Z0RBitaxVwSADTdErrKDlPkt8Huz3WPjyc5xhuP1575pno1K
b9UavSbjSnHVBKF8vbjzIenWTDXyQYAMVGy0FJsmt0cbGIqEb7FY2r4hLZ08yPEfl55KniSz2PdM
K+q4edwPDabNdLV6OpqEo7PEqc8v0hKSJTXPX6Xk+Sp3OA110weJgwqkp65GWjxUpTw6YkCNbX60
USJCRw7uUDC5hkXVng8UfaNIyIY85CISpQ36eprDz25c4c5PnQ3x7eYVnuyzlqqlYXLvy8N8zd7j
osDuMhEK3ZW8lyB8Rob4EEgcVOxSfihFtLIker3hJfaQpHZnlDmCpUyR1HUkDOK7Wksu9VK9T/o4
M6/TdoO+zrFtzmtx+aCZtRTUisK+VKn32Nyn1ldEn++2afxjex+flXUaP90X+On/yrv31IfG5yPf
/LAAwgvfC21PkMkKgFCEskDxkzmnoRifeFoqZeEr/FCHilYsoeT/mA7kVysKTFhRjfhehb5QHmD3
CDu/u32ZWTSgclT96MwHSX3DGfVuBapemCAYOCTQ1TZN2mzA0BPPsy77Iw+eBxZxU6PkGmlH87dD
zYY5iRwELHnC29HcjliHeptZOq3T3sLIvRrodW/Mz5dek0H+7Cr9GPhGTnCcO1V0WeQ4go0O1mEM
JnMPgAJmQJVuw6AAqsKQoRSOkQQghYUD/CqdFcXKxlu9YkUWmgro433I66ClVfuQ65I5D2S4uDGI
T+newdSFTr7+GO2eHSQThFmq+vYDERowFw6j7MQowJEiRPaeqfKMdd6YSyNvF9gCDeGMnwLgEKHO
ee1xnA6Q0J7G2h7SW89MdhcPVCz8aLXAgAl0HwMOH1zrrFzb976kGlWiaI1KrWChMfgmlYZ7E1GL
rdwr3mJ5dLpbLmUG7mhxL1ojp+W4TJIN0/HdYu7oxO1/iFe/WL+JQj+ltAPV4fsEh4//IY3aML2r
yxXf/swkppo4xAF3cr+Kr2fOs2qKC9qdh9z09q3oUjuQ0W4J0pwoKVIVYrbSDmpDlyrQIxIg5lS3
SQDKmG0uULyg6Cp4ykkKpumLiQMV3GFWCNDKMneowtyDcRyOoltaZWmEcP2wP/DFmj5S+QYv64Iw
nDyFNWIj0FRM9FNT6v/qEK5nIOdYw0Yt8lZvPE1LxjeAzq0E0Bz8kb0O8iajgnA4vMnLlR3SRBdk
noKtb8HRCyvYfn0SFcxwVL5b/5dyIALayRhDt2FfiEnC3fc2r9Njh1fdwqXXG2RAd0UQFfuViPXr
IA9rVgDEn4gaaENwIPE0LeIBvTXhjm8Cbw89UvKuIWydKkeMyNK3EgxcUQQ8sm+MZ1t7iC0u6qcI
WdH55gAsqumciiouSI5wXAh9ynfnkdK6cM4gxoRlKpFgJg0KnPlqlN7jzWw/l9RrWqoJNmEAeH25
7llNLdeEQledGQpVxx2iFmjZ+2CRIhVG0KvngCK3b6JZptqLoEKmoH4GxFBJu+gzbaYml/lnzZbN
WGotM7mGA+vFGWbV0uk3NGdYrVn5wJB/vUSjvEqsI6PbqCUu4nPHnAIkzvP3XAeuukiVTEjbNEkM
Sfo6rI+NRc+X+axY+skYsrxufMR/SV8TKKH90IJLcVeWUhadRACotdrksyHHyJ1bxK/iOkS9gCBC
IRNbrxKit4BmcHSqNlKqO4M1q2UzDDNT9t5GHVIf8NLIW2kChbNcckCGaYeMtEuYC3onx9SssFT8
WXWz0Egy2IywA9N34aIjz/c4Ii4wkjHpe35r6F6m6+6KC/e3N7ssknO5dX50AXTXhtYw5S+F7UsS
fIP4u4bRVBYlsOT5pVMJZgJs1YbT0muc+6GqBO5z55mnRd2qHW0hPp07X/S6ZbWRtH9idMlPolZO
NoG/M8IakRZCYbfdGgxHLQYhXdi4TDoR3o/lcTNZwvcfO2CKxoxTqTff1FJD7aky+Bksibbq52vD
tl7eK28C8MEvA93Tc35dp0GfLmAAoWEEU0L7bgSitA60xRjrnWZe6gZslim9FLffOyxLvn8JBqVL
6mWko5xQTvGO4txatQDiWSI8S+eYzoPXCWB8WfSM/mPzCQ4FB6oMrHD30uCk1c2kL+Dk9ugLCuNT
gI62cwW/cKJKeiAZKoTjNn03Eoql40knP9dYqPbcghg8x72yQcYntUCSLJwTEM86nwoY43hH2GHC
OjTCyKZXp4AnRkl5F5NIL7b6MX6S6PNZXmjSMgqJDLSH1OlhBSeZ72m0hZAQc9l0UtH5+SEsgLEK
l7PKKZwRZIOHOxA+leHizMh8jfhPd8OaZGY42GMNJmzHDyUEdppHfcrsZsrZZqhnPoNd8kiKka5K
h2d4p/gK6csg3OdEm1RfDcnJLW1lSi0pl30BZXkBsDCkCLTmi8uK+mlQkLuOOnVdndISo+Fs9dE6
TjpDyUXJ2J/Pakvj0dPGfCXeGutQJTZ/+pAoVAEd3iLZydSSy8VZ3UMiWt4k/8R5vteB0Ea9UZtC
sPv/b2FhmTB2bE5bJbe9TVB8LNi74Qb9AgGbYWc3CAL4pWDH4i8TfJO5ta7iQu+38quyhVsX4Dn0
BeEL96+fFAQv+nSOUn8FNt2jccHkOz9l56grLaHRH08fbNZJ5Mf8nAuJ5Lsz4gsFmCLesi0pLmbC
YaXGKOPVEAQaVGk45UMgHuuEnoo8xtlocMiAXFLe3sK7bmA907fys0rWcYEBSngjO+aXb2Q3WzWN
pxOu52U0Uuxq54CZcTMCqLQKuHe7Kjut9n4LmZwnA3jrD1pMkXjqe6sfFo87NLcqlzItT1QStz7u
NTiObZYBS5L9T/lAe6IxyKR+HX7dFAb3+ed7mIAXelcBq6lfOEuZNEYZhG7BCLmOA+aZJNQOFPz4
GZqLuBME88Ht847AQvBJZyUXTp/czkaV/eqUeMQY8lOyoJef2bgqFdg/7VOp/T+fgTTRf9MJKLeh
hhT47ogX5kj4WirD6LTOnida0imWc8DZgK9ElxBVbgF0La0kEvz+qX7PP2f4AWKNIC8Ii7FwdGv8
20fQGSZFn72Djvjx4edFBL/PaA0Xzr3NUPjUbADBwlyLOAKYiRWVDyuxwZTOeatpSIF0DlGOHHCB
36l5yAk5bhujxWTkBbBOfsJEten6/Zth9fj0W0sUvWYI4ZthawQlitX97Z2WJzjir6p+9znljUXq
V3uyaOae6RZoFHUTdRBbf1ECrMjqVlpb6W8ghSQUOcYw+4xPOcH6culp7W4kxQUOj7iaJ+0uKGYJ
+XPXIqUjdPznBtqHZlkdPW+4JgFtWpAPioH9wF/8zMrl4/zD2i6D4tq/L/5LUmiaTYVeLlldiTQT
x/bm0IH/qv7fvh5j6tjpkp5O5TbJpIS37mGuNyhJ4EaniYKvFc/WomCJQWVB4yleDFM4db7FUeVd
YBW3SAY2tTyIbRslThkSHRYA51dVZNDWAxu4F7NUBU3dcCrvqkli+PiFgkxzjwf3BEEO31ZM6uPw
njiCqW580Afz8T/D2heVlvyAc+tY0xhjjeHZcAwGn6+pBovj5PL8rF/9m2gjGzlJKH7HgA04IwSq
iyPAaDq2jvqfFQALO9ISNXQ7/ImcMPmanzKv7P2xGZdzFhj/9UlG1XglQzxhrD8gL4XjNR1/IExo
Lqbd/tpAoxg3HJs+EgRvKf5rTwokOFq9v2Vb7J2QFp3Egi+1LEQ/iF8QTuIyzHce0UGzYrjGePH0
UisofFGa6hwEFVeaPmzdxtgXTswjnia1UBxuumpjZEGBwp7cdF13bq4N8keiy+8kXz4rZfm41efm
1jeo0rUgIJHbO4XxGPGd7VLL5LRJch5UDi5RPmfvFPSfHB1BZD1G/v5wpG/jpTHcaLgjm6Ygf6QN
6TUjlB98OHug6qrYbxC+eG6v1HHhXiI5yslnFOhYQWKRo0gXPEQ/CJxXbaYXhz3Lt/y7CqREeEF/
IsARp/5VMgvymVMPx1UPb4IJdt3KL7p98HiZ9R2ZP8PaLF9DD8huz/BNzc5LZgPYiBKBOCU3sOS4
wyOj2RaB6Muw5luZYvccaOtyNMftpWsIOTbIvc+s0IgypIh7OT2+TmMexa3CPdLQgFsIBxjn8pTi
MR0kDKDa5ed08faX9RxfIRpvJRu//vLd+NqgLl8kIqt615A/qZE7vnobkf+4ukGBRKnMtIXj0wLz
k60GNFs1uQHa3ivuk8rSg/wetMX3IXGzfy6zOohIayPFzWK+E8n+Y8oaODj6K8GSNIJ+37Wk/Vwr
pMpRfPn8SgeMLYjJedR+iHVRMBygMowfOJvB670gq2SgUOOqpCNnZlkfJQQ0E+DiSYEPDvKjUskY
r6kM8PUltsdvZ4t5+Bdr5DL/K2cR4XaHo697om9iN3m+ZqQwxO8L/QcaRz0varcJw+IssPAtlWS/
poADX/gFRdN1VnSMDkGyRvdzr3euKwqj+wSFw+V8FdSH0qXsfJQgtsPAfitdw9fbYvyJOzRrO/zo
WsffyFLH0PA9MnHm7rTQ9TSC879qNZrPpOBE2euBNSwgbIScvGom/x+3RM5PlFwCRmTcmxDDW7RN
78IsflHS3IrOcU1Zonm4E6umoC5CcBbr5gdT4djwwm3DGteCa06Liz9kP33pwKaDiSkPnlexpfxl
XwsvqJWAs1TzwxYx8ENp8ipngM8TUpBE0iwNQVD2fgGEDn4QKLB9lvpDeGL1goO67WCcUb2Ttsq1
CrDvdzzlfDv4EFQd7liPS22XtKnnFV0LYY2/R6K1+aFki3pp9oFezZtacLwFCUc50722rlNeIc14
M+Nb+scl3t1YK+fQiQBNjNsZ9a4bVhbC7iFqNfRmp2pXS44MDwPfx3Q5iHeAqCcCmznarS6zpDI2
En5EhLWJne3RvEupg/nKA3UOcmrmVPn/Pd128nYJaWJOpJ1R6xlqoSaENXqDZ7N8rXsEPGUuXV5K
ry28RkrxYCzodYi3gPzD8+fZW+nAF/c+VYgQx0JbRNBK1zALsuW/wTkTTh/4qovvvhDX3IcQPC2L
P4NT+XKr+r8c7g8/nrgI1BWl1QUVSJ3n4hIezqXWRxuxWXiDAFLAyW36Vb/QyD6bHXFcDxiS6Ozc
Ev8C4dDdDMjCLgF79yu/hz+Cm2JHZF5laqoSR+umTnP9kPEBI1MxZjn8GTSlJPSO/JzLktbOcKvN
DfmnYAnv6CEBzcgCbDLgzBwNsr6Td9NHlBIJ3OlueryOV/FRjAu+E+qOyJOicK5wO9OjEc/+FWug
0vn+9rvQ9dUWDk6AoKw9pjrRSuEr98l4vOgZaWZF7HPTach8vcSr8M/1BwZLWKHxloms3KeR7wmE
uHNWnkhFtJ/qcuD0/uSY6EXmaG1xWzj+rOqoEBzN3UgSD3A12oIqKy6ndNaGagkpcvT3vBH7UMv5
pJd0yntds27msjIG+m+QhSHl/3beyq9vTSmzKQtDcyGxBWH8xMPH9RT+9Z8TmWlPucFgrj/zgvnW
Bi8FXi2LZW1DK+czKiI/xF9803wcWxgDHs20B/Kf5+/3Yp0Yx01t95w9WuCvtQo5xwcRo0Xk0BvN
kuwbtkYE+GjvACutRlzWI1hQ3I/udFgSD6wvC4ko9sa6xNECshnvhSnd8sRYG5mMtAZGXKiGI0ru
LA+bMWPScNtNUfKSjpfQdl1HkQDZ8Qs5c0uyRF+DXLVeGRmjoMKW/Q3FZSwxsC9lJMqvAOIgvRPD
+mAQQpG+ucyoH3mOo7Xz5qGwm/S4lhy0sLvX71pnquPY6BQOpUXjGyKr6QbcCHoPTdSRoNvJFJYR
QsJygU4yc9UdArHzSxoNvT7/bx8cdyFLx/RiBlVOtV1Ntl7WGw4ovZpoK5Y90P7Vh64Zbtm80UVQ
wLdx/tk4355CNZoie6KpuhOtJf6BMv1GGETGv76UWnuWjfRf3ZOY3rHT6tXcL4xwMTaYqcCo7SKv
Y3NZc0OtigEtF1IwQ6nc8FMU3JJ3Sw2Hnls3oCCOE8MIfbcL2j0uKQzOTrJd31aTLqNyFalq9lAz
5I0jR7sBIYqip3lJmFe/CusvseXGcc+OTUXMQ3UZjL0Nc97OjkDc6c+Z4YlPshgKXgLNtoC3rD91
+bDYbReqkci1lZ3m1PLWDWVXl2amSg5TACC/ykf8TxZrjCgeyisIUulY+h+lawEnOieICdY4anem
9+sdmFQj90YVO3rGNqrQDeTKNrgpgarGuG95WoNEyW8iACoNCvDbe23PoorGvB3q8LAfhAafbWoq
2az7g7F72NNpK/elciwrq0CqV6zdmGeWufoR5v7lezV3juHZbLB/Um5IvP6bC+RV+Y+T0paLhAIV
Iq9ITAXCDstDgcIsGTFPI5QEKuGNAywSFFFS6L/L5NRpZxUL6lHEZpARWERq14nGHUo2t05JqsCT
A3Q8jTkAoyKzD1ac2eTmO55sYMgI2tCP7/H1tiJ7n0a/+1bglSej4ilp44zb5oBe4iQJ2KwIjExY
rSTII2UONrd0PN5K9AkJnkUQ7Uteo4x+O6PU+wP977sMSoF+Rr3rqC3Y03Xgnky4EvKpp0W3rMi8
ihs4p1tFIg/olcHLMziBXqOIY4HUgyz3Z+Eqpj5yb6ahoc2UNcVXxBkNEktkdKQ5LWJMyfkOakOi
K/Yc8WqA6h8/R204iR8j8c0MqbyEtRykPEnDca90LpS0JkDjXkfg5QokuQBNrAOzmLGo1wOg/3B+
kRcQZQYHsnnYDKE6b7/svSkyFpm5xNmpQkEJBzNoKEtNKKJzZb0WJ7zUek9hsAdpCEC+k4NyNXo4
mMZ8dCxXvZna4+yTvwhGxos0lV7MTCR0ufqEA04WRkkWtSJzihLfYTAiiauArzU8020YzzFJW6V/
vIyXGD6eRIPRKtpT3oTNobC4zfARi2RUq9ul0SYJKFmtyAyqKJqzQNtCAhrMnp8FEuhzKYnIs/cR
IXqZJ1ankKtLRe1uRSB/0tbQYUaElQWSqxVjbv2F3WCaDQSLwK6zn+pwX+qxXll79mYk/+X9gBXT
CtClnC9u/9kzW0hlPp0YMcoHlIropTHdCY1tvdzg8ZPzB1N2OdzQe/IqA7wNpnOnHtdpoa/JThIm
6v+PiHz+t2BJaTF4PHg46gWsPmB+ZFOLzA3WmSpSmS81BO92GEkQ6ZBJYzXoyTG2099fp6hGVUfI
w9pBCuXKftlaOWy7RrX6yxY60kyejlBlVKS9PZTKY5BRLNQyO2dr8nh5TktJiNtiLSRFiYkiVnIG
C4Gd+kDb1D9ssCJ4i+JgT7VjyQ2bGCULmJYBkdtbNyQiuWg6XmlhquSH9/vU5FK8ncV+QgeBZXiw
VzrsoLxwEov83f3toIbLziilQEfbz4Xms9IK4f8Go/gpKUd+jwNl+rkVJR0dNKyd5Qyaytrh19bg
oWEydcYVADlbENmTZBMcVyu3hAVF6c5nJVrTiuGAF2WWzFp/panSTP27+dyIrv4FSf68cJy2ZfwM
RB4c1LXfI7D3XFbnipXj+k13NQQFBYqbncqEAk0Fs6QqJtJq/83nA+ogBlgfgQEOAWMKaqZCXTIx
7QnUiKQ2Z0XXacIymybcQT6hMA+z9TErwUuZIpmP+2ANOH9o611pm1rNewoSFTpt/u912gJlIEqb
yNzSSfVusuyuMjl8xJZN2wwTg6+wNCXI4hzPt0W19J048hA+ytVJ43SA0cRpKW2JQsCRYZA9v1rm
wMOVt3EhsrHnbI3rT+Iz/fVkdtW6wx3OIbPVhkDHMSknurlaNVLqGWit/WnYK5B4+jBx8+k1LQMF
203OzjAti5n+2puDMuT68rfWHgKGV9qK4itDwjruaj3+sztYIhrmpTr+9tqhAVizyUvrAT6qIIja
erXyVzuFOm9j2oRXAQFYY7bVpVIeTCBnvyceyBhOw/H2W5PjA5pq0+ydvzIbYEnemnKsS9+pAksT
Fr5pi8oof5fZhpoXROPLg0L7gvBxz0ICGbu8UuyVSWT43L4cDd5BSvHbKyg537KiuOyWA5v6VQTa
899WGCNuaFPTyaZFgswx6xS45kk9yU/lwOzEGE474t1iJlT+Vt+BHcmFnnnAvX6yypc8MdYlrsqa
V588HTKgY/C3eidfDe+iZ7us8NBphZMbWW9H433A9Dga4/kgagpaKKdJ30xg6V9U+wzICcpkjos1
9wtdF5kpxJjzaBr2lJEEsxdY93mXsK4E5k0gUxGtNDcylTuLP6xEF3UvQW/MiaJ4kyWDW9TPQVJW
2BmZoqlL8PC3c4e4Y03V57ADj96WAycopzb+Xfr/jNYhab0jloNLzcfXqhcTQ4zOALsHp+4to7OO
HWKhg5ShutScPtoqFk4nNnV5pKRKRQ1eQojB3LKnSHkYDfXDL98J7Mg9U7k07r86pBGQNrMNjdVc
2UyiDt3R7ph4+18F6mqa9foxDklbA6TA/QKsdA5i7dPeUSogX3f4iTmSqETyE7QDz+lXLUO2DBAl
LLuEIkAPlEsubBHRuf0lUPEjDa6aaXPQ6Ei5irR0DW0Sqpdgn2yMIOEhVbODLeU4RLiDaoAVH4b3
lC1Da+GpU0rVKEnkGb+Y+uTSbxlclS+TrlznGb0hyWFlzn50vzDfZSmGEyole7DYLuW3IWAH/5MZ
1LzLCmBBHnicaMQHAwu7DpLOmSBxrN0elv5mSk1Ge6xMApClHyAY5LH2lx9PglBhyD7U94BCxcPW
R4oZtX5t+T76cAtmH5cI/n7LhNuYRj1d1TKr0WWdSEa8fkIQQyTA6IoC1XzhaKcmpw97xJkgMf/T
vlU0YF8S06OfwndFnRx1KsjCIbnDn6mb8wu1VMn25o5CclsBy0rJ4GHtBbdSgPbZhTWMjJCytO0s
UuNlx4g9DUay2ZvNV8+BcIcXf+1vR0OFKPRSV+ne2/AL955NkENPc6VHctiUEsV+hB0Es43isMN0
fr/r2G/wpw0DBYHHCozhNwoCzy9aM7AxuQ6zNPjOqzlxwXTf2/M6U5QWMoWh4NmKJZ0bfI9ShkKi
OxyZO1onRFJ3AWFBqpfRdGgrNxyRBFjJhB9tl5MELZVbNKIs/imMksfPe6kUIDJzGyMU0w/cAU0I
bvdiRugMm6hzl1LCvgiJjeFO63CEyPQpkZz4dCikfWgAL9zJ26DHDilsHX0YhwYPw1Q6N/jk2ep/
it//vt5u/PltEOW/y4o057OGixCusx/TNecz0ocn9ZEz9z28yIUjL9vbccQHn3V40NxpLTK3pC1c
F5dEOBCxTxCtTdD+dJm0u9Ng0hXwdCd2LM/DWZr0i85Nxzh+/Eaba/+4ZzqFi/0m8NRqliVDMcvu
At8+yqJk089WsClc8gIyjPHFe/oY6uesxk1rnJj4VOg2xIaH9vN2ZgzmPMKHee2IEMCl6cSp4UfQ
0+eRX5l1WvzzNCoPncBjH5aI3laAcrfDr4J7OG827pt8rtna7GCNF+J43aHiKSBiIYlIMTsTNcvQ
PQbvxIT0xgwQszmAjJHUfv7+q9UN1wxCqro508XTGfF1bAcaEpvlrYWhRGe3Dd14t/7uA2vBWxWj
5Rk4MuF+96W6FTFNtkejwRchktINPsJwkptEMilYGJXl/YSgIGi3Xm7e+VXx+j01hBpGbyAQ1F2K
CABd194p933fKfRXbYbUxGPho0mO0TPGs/NRtUS2kFYFt/mIHU1rrQUec09k9mdeU9X8NTTbHJUx
HqtLAghaooxtNq5f9vT7/+fRgxMH75nauTGiKGubcUBY5d1255tzqYwaUO3utlpQH26g13zt/HzX
cIoI5+EVTsp/k6m1653ifLN6ToU86ESy3mgX1yucuB7z2mQyOu3PnMiTuuM3FcctiH39VYUBEtDi
FLp9cHk8ll+Z+KkAyKTItJtChq7/lkmCbwng+uBkUNIIvEKVQGJUCE/BlAePKqnDPAdnjCuUftIs
ht9yHLX1SwvoIK+ORt8mcwxO6yNoeIyFMnm6qDH20Ei92+EFXMK7Z+q/hTwuqHRwVFZWDIFAZa0j
xnvETIA95Qbzll2qLSN+JeT5ev1dYW8ndDtTiVMF5FNTmvXRJlN1emL6TXFqdZwihEHkgUA6glAK
ZhNsE0BqYkTxRAt8vEaXj+CYmEeJXUK77E3J74WsmPROZLJE5P2wv1K6VNXfBIxIBiDjCHV9ItXX
pDiv7YJrQFD5TnpFPZPey5nIpLSsXcS8WL1CPCgOW+D97NtnDH+Cv836t74q4aZbTgu7FmyFS7pa
1hrep7dEOw5/wqpj7qIUeaGhSlDnwBVU3ovHSvwU8FIl3huxofO2Ikt92eE994VOuJConeIBI0sc
dgqYpD4IK8Wp+PyHAFzXHs688lsDfat3naOn569TeNN9LF3ym0NAr5JXv5+Br9SJh3oKdTDox+bW
pyyzXfpitSybw34wiSLalWJfBlNKUQQVBo+/3TXBBuc2DjJXhMkL9X1AyYelFQJsxn4xt8GgdOBo
y9IpshcZDq7M9mWdiicwkz4687v9gL/+kqyJM1s7qTgSn4sXnsZhww4kS605miVtlUAaiJAlznoa
zsC1uUGTsArkCcldzIHGw458Jxq8qD7+/1HFiwAQksAl1omMRNDCXqTX/B6YTEv9ay9Wsb3D44xU
7lyqruKuVmqLvVQm96iNWvCI4woaWsxY+jwo4qjwsHfHJBKeTXmUStJImkCvs72r4L/DPC36mffp
Qw8Z7mhf4FG0hrUJpyl5fG256k2ZKJZeyqoCPjchSuAHN31L+NlYxqcyGQ2mATcNqnCnP0ck3Mfx
3rvzvpGzBohpM/G+LJTQsFVs8+aVWdRxFUG+Wr2C4oKKONpGrrcvJ7iMxIq4OD6hals3kk1rS7QE
35Ak++aS8EviWCdziPXAFvt5cUfRVwQ0MOSSNnJRqFMJOySFgA1KErg3pBmKf7P0UaDdLnbcf4fa
a8pAPu68Z9wYqi3/AQkMwz3KWEcyQyiVNcDBEEVul3b3sX5v8z3sceDnLqFM9OXLYUYd3zR5f0MH
ZJyt2wB7VJiM/Xahe9xaVwCeFnpDGhUPrxjD/3qJD26yC5CH7bWB3J9OKWRZcyc8AKrSSjJGBsFp
yacXgp04JpPab8xFRVAOudtYkqi2wLmXRzg01jhNPK4YsM2Q/zsQocatyEBPjLdSRtVqaXhpwdrD
Z4c7vSxDKwHN3SUsEtFevGEXSXaG5Pw0b86aVIvNLqYTy6KKuka9mOrN7KQnupswauj4WrIzSbu9
3jI4GV616fI7LyxRpy9XA9CtjwUccj++mRKdSqWOAWfMo6Jnch2HFGLk+UHDiI+Po6bqHbRbO2yX
fjTWmaPxhEBuWtLgcjMctd2hrFuWTdX6NDtVUZpJVo+AQOPyaB2TTN+rOAZeo2o+Y65+VZu4J2x9
dXbZ6VSzqe++v3hCX5d9ugjbWVJY+ICkyKgMZXUYusiTOAC4XsDcgmmS5Qjy/1g+rtil3TpKOj0F
seV5VEkU0bghTpeXGr2jSD9vKyJwuSYx2MhPVcGleVxL/9RKXc6TU1GBj+SNRVow0jpTkQAhe5od
Ss2tGMTPWe9ZrOMoXuJJoTmsTNigD1F+fKY1vJe2NTySaK6hxT2SM5ZcGnf6aMb+qlqPHx03qBLt
GzHITtKIe5gBkrC2zydC1JsQ/5tv4qouc1FZvVRGWMGOrRG0823k2FX6DRLawmZdXpMbCIrBpPoR
LaVn8Zd0Tg6HjurPV0RJTvh4jy5vA04LnsHZKE8/BUz6sonhEPBDzkUu7PVwCAK70V/H3YATbyYv
lK0hTL8S3JHYsHbNb1cqQhxQ24GWEfwzrikeg/PPFfh/2fLsqsWRJy621Q1MKx3yyAVBGf9NtwNw
WuhxEemGD7M1LVAV/cVBSdtbIZnjosmJmI9DqwYk/rCzDV0RCCh2rIawoGTD05WH56AUS9K1FbrF
lgzzhnOoGHszkj0xbZUXFmsASeWvXOmeZ5BKZpr/OP1mwrZObowBVUEPGS9hNbD4O3Yy+9a8ptci
YqZjOsI+igmC5bo70lcY5qyyuREyLDO5WRu5Es8frOM8/NyiNLSvpE6rANg5DI6TY5B1aq0VXs7c
HkWDKZaqch3+NQkw1jEE9xGOE7v88lNHBxLFnQf/bNovoLVj5N12fKu1AMPUqkKa/5bIG6JreR24
3+frFRUJxvv3NmT2Tgi4ycKNk4jmsimPe4tEzjJfd6LVHH2LZH1rm0FuRdW8C5/HSxbGXg3APNx0
kH0hySt9m/bm1fp7SGfbvMLO9UIz+jCbQiw4bcdX/oqumcwK0JzITAJFPdh/cTugLidd+2E8x/wr
rEwwrcOnlFcScLbNCnJmF8LzAMsuQ2cFPUiX8icYJfD5BVkn0t8RllDkPAgim5EJvvnwWGpJmo2q
xHQ1xwHcS9XLeJUURlRF81nzix7bagkd/DsrnT8IC1S5d2i4b7DAHbEwsN+YNASnUVpVBozfa2+o
ZGznQYrfmza99laKdpmJFVX7O5c8lg7sOZ7zOhfkFfBCat3C9WJWIKRQvYKhEbK2gy9pQVKpwuaV
y0CqgobmopQ/dQKySPPh0yL90wAej12RQGkWl9OAEvWpnlugOCX+0+bL1WpiCqAKWFB4oj1+oviJ
cCkQo97qxOvm67oyeN49sPqpj9m/Bjf4EJJKEKAymnPW/Sm5njNtVqlyWNsXFok+WHRLEHYwRp6l
JdeOOUASmujVPWUeaMsHIXJi+cVMGT83mOzLAVVyD5q6OCgEO1gGa1QKbWj1U265tO94fBUhp7zB
SgdJ51TQba1iACyWKqukR2RSonxvuqnzUncDYNI4J4omMPGgrPIg/P72TnS4brVPnj53Yl8eP7lO
zeZOuutV7A4VNZjleNrpLcw36CGfuLORuj+B01UjkRfemXF96y9vtD2m6Ei3LYlngv91RO9tF8FM
H3gP/Lud/Qz22la1wmp0kLF//0Ep2BnfK4JigCofYvBxGSvHd/FwTvW3pui+SnCefEYxdcSt70tm
cTt/uFzXcLuw5qFlNQFhHLzb2VotPOX4IIs0a3/+5k491WfAZTuqigBPVI7ucQj9iNmdRoyV6Hcg
t0ph6KMcgTfoLmruPMHpozq5Pyq/v69Ze/TxLDg8lq1ZtWRZz6r+rKdMTGhBUK3RuTTrvwThdGQa
E9wGekFe5DawQbeQBaQC9pSaDq1jWYcvIez4KH4nUTyd029lW5G0vfOIGvUE5mnWA3WsniCjFh0s
nWYKF/6uGb6KNXu7VK+3EdrqE5GvIZtlQ1yZ0YvpMttlSQJzQ9gMpfupAXYVHcMpK/aBSyYeSr8N
adiVbKP1mY44hxJLXgsB4oU0JVklCyfwDPba959AfTv7ujHQo/N/mwZ3n1EwzpMnHjrzcps8mMOO
4XnIC6YYFmwOh1983vZxHT5LPuUr0bHc8BUKmiyEgI+Fb8QYXlrQXz/5BQlK+phvGv+R8AT9n55i
TSHFgrYKez7WKjA0pqEx1qbEs+b00xeFWJvlI1v5/AnA90WROOw7AYnC/VHK0rPStQlJT3BXwOo8
fAwrr6QERbtrARZPN30OeA8Ot1JEKDDzHSZhrVjdMZmoC9n0Xv7pyESiek8VLECapxSsSbBGNYSH
J1GvTAT85s0flbaK3x2hnuHCTDp1C247M2UfM0JxLUDs/35scmav8sKfnsP1mk2WHZzBk4wg56eO
nYBvP/Mk5gkWoXzdVNv31CWg8/jF+kVUK8SUGL9mKQ00S3sZ86aaiOdaBejZgr3gSgyEt6NyKmC/
s5dukd1k4obRmLQM+Q6cFedKHm5nnqjus2kUozr8/G3+3615aKD68UbbUDCLr9F+Q1uLvHSgkLSq
h08pOtNRZ9mMnWxYubsOZhTMARo41cGlQJe8oYZVImshgDrzqDbcAR2jngzOHs8TZEkVvfHWBAGm
2lrm781Ndgj4v+FZ7dLLAVy1FbWl/6I2kCbDz5Z1trUSiAburqcMy16LQw0pJVAXLKcrf/IwyIIq
YypWy542rW44XT+XfN0M7sohW7yK+HIYh55Io3Kft6X4WrzcVsgKhTImjpNhYG/1pfMXvuDSoILG
jXTDsDpHzby49Nt7oXq91q864QuHfkiua55LdVwAx9PxfgPPay96umCt6uUDqkRWq6Too9WcQ2d7
m2hNKn+aqa8oxokUrc+87yF+cFkjQf8WdWlvgO/Cq8d1C0K99usyfolb0Ab9w9ZegBIwh9NrZuVM
Ss69Y69WfE6tsSslYzq0SBnj6gxGvlxTxyevAkOX+hLRPI00u5xEBt/8NkvnrMAO4L7XBQiBbrUw
egPHay7C071aCBSt6YEzVpftwBhzytXhFm2VdYr39212tHhwfgcMaWuorVPLm/HjIxqPG1WCQDYi
M47gbRzWyWmWS8DlE9bszLFQ0MiTF2jq3T6gqqiLi1XtnqRoDCWpTGyrYbyNlOhhJ/n4zMx2hTdH
6ehdfI19YbHEIUPdWqvXxyBmoewxu/EL8hFqgs60r1FB1sIT8BE3HCLEb3XDxzGUjnEjpbp1IdrA
GDzgeT3ccdOQObosX5av1xtEuVU7XQuIei72iN69GN+/+OXfF2UP8tx0jRj5UeVgyF83x9arf5LO
/4DF2krCE5eWSN3sX7gNtC+sHJ43hAPhZO/hE2fFMCnJ3UUJHC1WoRjV0CAJorniKyEZx4jiCh7t
baNHk/Zy/H8I/UkYQk3aHMu1AFk/QrZyoxhgGR+TeR6NEnlbbbyyxrXloL8K6eYrsoI4SQVDFmnl
usuefL3HDm2tlW9jK1g1FdUixpeloowKzsGbKmeWlxoBouxPFjCyxq8r8ODryTt38nIFkgqoKeVU
Uq0+bo1GhVZNJvkT79GsS8ViCyJzuCa70GGfZ5DmL1jDnpdRZph3Fo2BFWyVOZxTO6dh0uoWjrdL
FEjBfVcTCcJ+/rXLijDH+K0GIoUjEP3lPBiaCwpfKW/tr71U/s1k+NBbLanIJxA/y96oq4czzt6n
Klghtx8qwGsGh6If8zZNYEs+8advUizdEwMP1mVKq0s0iHUJBGSdFhnaeY2x1nL07Xd410vwe7Aw
R/YghfPpN/aFurZGwolzPAw5LI1Gn25ZldN5D70aVbnyXVLZHzflAnZY2PcbpF3EBWZbpb3OARZG
k7f+BlxukaStgm4Hn+NK2G2axltVekw7+GJwj2px7vt1m3ZhQgoLZ9FoewgNC8Kq0irZf2EtTSpa
dCfOVITdzgmF1tKln+LQlMIPSvyHPZOvT1AwAoopp6mmQHytg69CDIn310/NvVYAWjAb/K0t2GxD
EeGSHfF9XOnajkxPl2OTCyRg2D8eUGkqmp+EmbUyEoxYWFSd4HVG1vex/S49gFvOlpF70SGzjJhm
yHiUQWNhnENGZLGvPwArh4e+49ghh4WtkeIJbq9Z4dcfmb3oE5+0AjFZnTXPbVeHwWM1aEdlzsR1
xA7fJkySZ5xUiTx6K1U5HywkX8lPatt2C2gRCN9IE9VzhLKn0qLvIcaSY5LSRDb2EF8mibYnTGXw
M1jXK7ngbrwhCN7biUDnplaG6dBwPYjiNlNc8jbr1dy4+VH3AIvc4o68go8XhvIwqpAyxPUnGA33
9nd7V5jgNOvw8wmpH2JZUxWw5cMGzNlaqFR/8lmS+5Ie9JN7YXY3XimcsBzxSmRCbrz2iZd+AgYo
hV9+P5RsDXbfGjNalsigbyG9A1IEqQwHirIL8cp/Z+b2suIema+DLD7o8xT/CgkRHtVn78AZFkmK
6vgjv6f1KwjkArUSb/jCvfwnWSK+yvdhuI4boVEoXyQ+2YdLMC5WlwmyBsTDheFpEePwoGqQNhZb
7D4T8DjculgO/mnr61LeSLrsjf6Cd1EPp+TVE0C+/kUxYlVOF0AiqPP4SD4sd2aVA5OWrMQD+Zn6
MUMg+E6TeLyskRZlhuq2ha12K+2/Y9ms6mMlArYW6Xx4DiHvKagEtybl4ij1XWr+oq7sj8uLxcrW
bG9NHwUwQT4HIEAUYLlALrACTnqDG/x5OonjrWDKzmz3gWQZO1BmvVk9b7eWSA/CWIsS21Tqh2qc
L4m2fd39X9ojC7dhdfPWuDNnbLMELlSPDh6vfY8ficF3KHyv2MuVNGriOR5N7fKOpn03RW+ZC5ew
GL3nWoMSBZD7ytXNwl4M5RKyQV1mIuDS4UINaA1RZiJaUP5f0eJh6LwPFFtHsAsz6Bd7/GYMBMO2
J21vsbGS37RKfEB/E8Mry1z+qcicXosldxjpsBsbFm8yPTnnDypt2bEiffBABk9TxsffpenkV9U/
9uMcGiLcyefvACuu4dI0lDSdApYw04Px+dknxOSrqamEyvY4/Ocb12J2eWTbnRQNARE4bn2ubXmD
qA5fyf4HvBOUYwD6fsFGthLrbRsJ8LgEbEDgPVR+Sfm6o+gXUxgCdiUysmaE0yjDIutdrrMv4Sef
3ZOlMcwtzzMK4mz+ekTax3vpAXQ4C1joSBIbBglKQfwuk0/QkmFbb4S67YvY5IJyPuuM+s8fb2mG
Gr/Y/Ztlm/2uKMrybakG466TZrLu4aOQJQ1cxKlJZmdZG30lNGCUuygV+vHqKMEIDqnWjSY7YVz+
G08HH9WTlHQXcjeO6+KxcpwgFuMhj6U2mrGj0fAABRdF5/Xb6AkWbAcvq6yRdNm6QchMe3A+dwqA
Df2oOf9DfG0dHGtaHRYswAuvV5QcQvDhHe7paj05cb1598yjANC6nObPo9gZgHsbZcz9s+ILi54v
/RK8xmnoj+HohtcvIfyIyzaFWcZYuDyaTjHYPCgOGbhAyDTLBPi/IGZwFbaLPlCHYq9RW/XBSaRv
5wR0krDLnN4B104WxZu0td18BKWyd1nFYA/RA+8LNgbCn7AK6Qma3B4jEFETZcNo85HfeCp/fM0M
OEeYAOLhmgPDLH+/hnoXmF0KlD9LrTSWuB5o7R9aiWSq1cQ09pb4eyQDFlJd79XGRvTjGLZmd+xH
+bn4BRaXe088P1s/iThAy0lzF2jkLbNl40yh479wG0pnxwbcMiuED29fmUz+TxS6lRpzaMAgyqAL
98hcF8iknODEekBUTqV3/LDFmCCpySJbYNvzmOecWhrF5hD64ee9Lwc8n4ZEZwt0lqBPDfeb4RUZ
/OMP9PF4thmdhk14kyycAQqVzLr/UgwOI4rSocB5aIgzPT8LxmhCYlqmdxGZGZTMaQ6wNh+r+9YA
lloj/uULDShzTSjwNMXaVtgWw63a+jmd1GwSA5cmFLbCEdrFNoRX1EkOCH5BLarpjNAbpeVnV2rf
kngUva81c0VsEnY8vPCwjj/YFLSKDnENTnsPq/u1iNACjJ7FyHWDsHU5PnCv/fwyX9v9HOtc3djD
x+Ne2rQl8wnN0R6VgVmMstJwipO2wp9USsOlmdQ1tT13vwODYnPXiSLQSbzfcMPuRiQ2p78j/770
FY02uKiUSgT2CspKn02I8CP2JSPLWNZHy7fJNE9cFhpY7esdHELshK4f6Y8t214p4JhOT/Zf/Nvf
AXli0HOALAsOv66bd+MB49tvg+2O3uECHGY5hczjzN41l3y0WBJwSWV3zX647OphZpW7zsdns/Uj
/CtJmALH1CttDc28XBhu6z1zgVh3seF19pkKSxjk/7trI6W6jdgPrp5uU2fYIs9AM3I6G6eIgA2I
mz5XgJUvT6UWab2er0dFwgIPOyuGF6XY88LPR1pQuAfKFbalZhZlNlvxpz/S7m+mlYD6NEW+S6hh
Wmvf1gaevfvzeG8NmEvMferC1vHsVjZpAH0JdtboLktqZVHvMZ/5LPegUUG4NO3XGkdpy5p6fZxV
DRKtscic5TaPImBGkBb0ECx5anDpC/r5DbAk5mVP/eTPHLNgkNfu0CYS6L4v+xny/thfdqc73CPr
XzihH79wefsiEWapA5F/AK1G+OA5ZPEFiVYITfIMfzkoe8OFh8zy3yFlshYvdV5x/CovZnR55z0Y
bUC9yCafSwTnDv5f2diA8dAw9OVNI62KAi8XaokShEB/30HZLseXD97AQGPZ4Jy2/4XkXUZLHHlq
0mt678oDipBJ+G+AukUedL6Q8NOAqw2889tgNGI6YrtDFiShGIefeXPIwHfITBTLLLEvzOoz9F68
gYgRymLmPRC3mXhQzHDCXOZ+5lv4ScbzeR9XL/HApCqgwekTlxBwmx3EOk7O+zJ1z6S/N+7U6iQ6
bOBwhIKRXI8XEDdxpeyjOCMlBeot3AMagkfG3fV9qGVDyg2GnYlvKx+AVZxoYrPLY4Z0DhsDS7YZ
qVvU37yqB4JOf9Lu2zs69JvW+YW6ZCEA/F+dDzwjI8iFaU9USF/hkklP2PmclJQJ8YZaOuGviYah
SZLg5NpINOGbCYxQatif7rrVoeu3wYXSovHXXk38ldk5BMD2VxkjBbrBiVhCnz5UQhMp3KDWJp4v
3yTuQ+VyIQOFIeQo0mNKCcnxaYV4tllY704NheHk1Ohg2yDHbxgl/5ZZZPwJai2+d721ZhemMJPB
Xw9QAChv9tGRHB+ucItKbdCkz9W2SIHSaMeOr88W+YKKidNt4UWEi6avoP9pjXnZV6XV+sZlGpG3
26WZvNDBSc7779cxPBU6b9suWDR//P6++OwFz8xN3V0SufWGmnBVWQkvMqeSo4hI785pC1mIYejp
js1kDCE9j5qwrw6+qYFIi74Oq7j3ASAvGWG4UPgsXfw98VBnPCkvvPafJNZXtc7ED4h0mu5BT08g
rzsZPEipK27lAALZr5b8pLxabThn/TjCCGhSztD+stm5msS9cmih/5TKhXInXTrkRiLCrid9Q1us
JIXrlM4RzHnsmTwzI9hUJz5njrPpNiPNET3O3hR/JVjIqWCTp6F8CzvvQ0Oy/xJXIgIsKXmSKc6Y
xwDl0yJUqDEzRsIPu0SXCkwH1ssMcf0dzjeqhTha4FlszPNq8TzfKZHEq2OpyQwW46zPFWIwspbC
ONUkl7weOL+/pwe1YDUr9XlCA197kM5sC7NptkV8MH2OH8kGLipcPRZaEuBV1pjaldIjdLMUjJpo
nc/GqqqkUSLKOvfBEWPIik8SzDP2QksfsGHpL3yDC1ShJxqVgIBvW+KarfvLByOZ6YFBOvrkFSpw
A5KIgYzDwSYKiGFms8VCk1pHTXJkvB3FvZZa++ThLAd1vulxJpLNhFSbM4z3hrK9sm7dD286sks+
pTZxcTkz6lclWwdL2qDygNabVC5yq4XP5Xhzg0YJbPMT2J/Iy7vMVVo9PTeSfZlW6paEmf6LV6KX
8ipF7mO6B3J3iSPVRej3mL0VenHiweMli7faO1ZCP+PACH7RKbpRSs7MTM/flIMwLJ8Rbbxiw2S3
gBDhTR+BrWnanbRSQzPs4A/WsO4gjufMpmxQ4rVG3+XhM9Q4zHSa/i8nU3yh8+iTQCpxSdUQ1Ivp
3wK9Y7i7z+l2e5YrPOZE07UR1sZFF2Q/7ekHWgCuM1/Q8VlOjom7231XxM0C3QU+jz2btphuK35r
BhEFtQwPlEUU/PUIK6jLtmoibXT50v66DheqgWDWUJ81Gxx5YCCdE02UsaKcIMddwMujBcRjokNh
DWt1MfixhuDmBHt/FQdcisKt+eG5s1YyUaWjo0e7QOSTFOC5kb0javneGy8ht7ZJCTm0ujsruyDR
yOlp7wbY8lLbM7rTq4HVAQR+itQoZzus2qZSi6aaJffuWCQO+iNp1gly3ycLi5OvmuFgcnaUNyeJ
VBzUczp2zb/c5Oq7+MKIooX0bpZUGwbQg3HwaDcdw0vZwKjLSjWNpUvk/GSzFLW4S23O2u9MghZx
LrOb2m/Wm5gQCSeS1vQakhPVkw6AlGA79WEWM45CV47SyGfz+igsZEe/Js6as7gzAF2EnfvQL0mM
tkPDRn76qb4bliDJ07DNHeKMitmVKdadeQYPExCN50GQFQkiMkR2hPGcPAopIHBKyj+bqMMAauQn
xmm1pZzw8OmsrWIjxVXLw+AYmKmhMAOEPItcOhmppsUp4t3FZVTvaD5g+aTmrns7IysyE7yDNEJD
AVgJWZcnUo8XOCjADqVJ5WUBKdM91LouuFt1EFMD99SypIFkmr0sBof0Xxnfd7zmCXoril0ep/f+
MyMmKbjGd+EfEzZbol/LKZVDJaWqsZaPOZHX7zWxU28dQXuOD0tASPhhu4bnd4UH8DtW9IVfJD++
44O2JCRZ1dhVFcSgGAXPBrgH7YTUBtLHQ9SG4HG8Bl+UcKwPmNIuKlt+ay5D5KF/i3RWbe+uq3ed
8raUrpl//6yXF0WEC3yhQEOs7AwismSiOZhfqUOlPambBP5Vo+n4eLEjAR75iPxQSLSA6CKX7ezH
2X4eK5JYo4g7w+fkHIYjFNwUwNQWKu0mBSs1VC3uHbJPUMYq9i172NKee6Pc1N0/eSZkix9I9rR6
6P9lYbMngkLhgv1CwxjyDhFcXyzwb8NoEk4UYgCReQDM7kTG5XyIjw93cGtuEllSU5G4tuQc4VOI
62fsCTeiEq0qbj/N7HZNBy1FiN0yAL9rp44Ebxd1ntYd7Ga2FbNbWv3cu20OklNrz6IUY9JjQexP
I9bkMNd9bYR/oQEjD0ycKIX3BViNEQ/gSuHEVFGbye4d4jqYgGwVtyyQWcc4ES04mJhqaONlGGDt
kzBaWweVfsMT3s3ylnIbi9RZWbrRMWgc/wM5fC18BzcgX+NrkuYC57YMn7qYy2ayXXL2kRYnpoCc
QNZqDaLued+FRWbkEjnxrRaNCTFB9VDf07xtwwUsgBxblIq9aY3xrjaB4phyYxpi6dFEAHYW1JUi
Eq6gGQ7Dh1XPg/qBQm/SziWx/mdfK1goKkMN5K+dhBMuGCgUp0sOn8Ay/DfVkjbm1wy74z7FOMfc
438ikJWm5bARSBMIladbbHG69L7OwHsIYzwV8U4EWJ6uC6CkTOCHK1CjHPdGNTpz/xJdEqQ9OcGO
NtK6ih4Xz3g95xLea0iziVmR7OP70c5SnT45mD0hlL3ICtD1e886oBvNZovovoWM9YzjziSk1ZOG
ig8bfmRj2l/QhJSUy/tO97LRzRRj6t1ykyOlODQHOqlWkh5bUbnUHNOfpM+UwoA23hgQg8/1KPbZ
IdJGPAVRalLri9dv/AvG6c4xDi0rdsmNF/AiVXdAUy3fVcHPhKAt9O4dtTxwzGD/DFXA3IrXPxuc
54MGMDmfAEw2zMYJb+QOIrmaNRiHQZqVpYv2w6x7Th4GL3d9w3NpoywO+VrBgqbhRpcbwHxu/Ek0
TGbVafWZccnsTXS9lwVW4D2/bgfq5NyUXznCh+PWtPLjPUME4NpFL97pU0QCG5Q6/fTc76NQ9vpG
jJ5sIxBMDWoOHzRmdrvjqcV2q7D5XzSdxqRkk5PEILrxUzoU/yXrLF6cFD2FBfkefa7L5Y+Av7HC
DjIUj12yHh3L06BVIPgNDvca11YQxFi4l56YEU57kKiLqOJwUdsLrgfr/qYvvjIox4qm9w+UArZj
wSrf8BoBDNYE3M6lWYQgvQtyxNBPVy0usbiOaGVNkTB0TpqRqxgVzc/2QYif/bJqVWSw9CPPPzI/
EpMprviY3tOyhBUdM8jql2nwZssmTgw+SkRq1dFVoAdWkCQAQGZ/yCeYYIoc9JkArjwf9x83d0vj
M0MEUkHMNWvcImrPswfb/yRWWlukQUeyiHTs+LKDFKXzncN2oenF50nPY3fCQf5107inSwKOpZpQ
eFIGo+gLd6pPi9y0nRK0wOxEaOc0b/ShwZMw6DwYthUyMgdjokT6WY++HjPah4Y+Wn+dP9RTD+Q+
tbqlx6M5S7qV0CSSW5CvBXCw+ft2vg9GQotRR0YPGwJOgiwx3+NJluXmUOxKfsfZidAGTyiLWTGi
Xw7ZcIDHrK458TQakQDs+TPOLxNLJYVjXY6kguTEO2UhiaDMCgFh9UlNGkBy8feA7CfkSj10icBN
oaUJVs4D6N7nDLWieNGr6Jv7dY5QaMLi8SuUfl2nZQjZtUrZFWn3P/bfz3j0HD8vK3iYmiWoOL67
C3r7nffvShtXWX3waofQsg9cyU/Wv5z0AkMWMP1jvGbohL6hLxBPeNAUJHqz5FsDDkIHa+GmNZ8j
ZtiFln+F6UJoxpBEfBVfSo1xBzyd5OzCTAAA7b5TTrl+NZffbBZ0eTn0JH3E8kVz4zSXCQNkCVOe
FV86swqW29V2WgLvntAKjmMIstIt1wFNoS2AtFNX0QKf6whsyIcT1aK+OpphxxhON8iRZ+pAKIim
RUPpuscH9Iwc2eFN2osQW0BXZAeVZQB/jqtqwdeZYfGgVVg7oPfM49RYT4A8lbVD06nOLrChpTMH
4LsPDkP5+aIw1ypJumCIontGny7ozJD8itDd06kXiEzy4y3Bq87YDSsNzntyk9mXq5aokCOXnMAL
rdIaX2Kw0vqc6QJadk4A42ypOMJMn3s3a9cnpLQeSumLdRzeJ6PvUyRyVGChzwvg8JV28p1bws8b
v7lMIpbchw/97GrY60yxSdmklx5YwLAWKXsBwl8f0+jJ2btqL6Uvzn9dCSXtul0tn6op3J+pFZAO
0aOhgwv03pb0B6A+47BMG+tfuMWl0Q0ZjgzoKJOl5zQLDDnEE2uflSkeXEXck7yBoICZHyUzyv18
tvbUWjkbrRob+iAVACU6evuDvGT9CIR++D4hht67MLk1692/jsZUqnJuXwvPQp8DdUXKINIKU1Ib
AzDoZwghDdCPurbuuUeztc5iYJzfHoeHZrGFxLU4lMOjB+rnGWJuKHuHE8dqbrfx5A8aSB+xx5hp
dHERsg7F2y7EXh4n7QTPxYCWLAB9gJMOnCJKkzvB6RO/giX2ax4CYzSS8z+Tr+3R2bWjJdgtxrVv
6YqNnKYvPbMfn7fMYXaGjVTlNn+QrNinhvgFziOROr5JBkmU+hngQH2zSJzjkxBQq8lWv0CLNBqY
KYonOCjWexPh8iiLIx16mqh4lpwyk3yRjkU3NQols80kEujg4j8ZOBNJPeBd1Z1ElX07RB0QGW/g
+WzOR3Wa8RaRHpkbN1Su3KujAiXNaQ+LLPi6W3XY44G2dqGUoqwfKj8+autre0NsBD8o1WF5qpOw
4MNEON1X0M4jw0B+kNIIrhNUmXr5+2CRSQ1zNDqeS7ap0JEZfsIyE9tN0hUP7tZpcZr/Neqd9wiE
693nC/xElS48iOrmYL4I7VO+f7s8QV2ureY/PbI+mpniQlJsKvlSGwzo3J0c2WNBIySNsbfOkEgP
0m+WhSxr2eejq27DvDELfpIFrzpxyltaODrKTORgS5M8CjI8llzpIMOsKD67H26EBcEraZPmYYLY
N5TqbIGQ9sMKzBACt06dmHbLkobeqsIAN1h9bssRHjq5P9s4vH/KIRGA2hQJXw0WvfslZvBFkNP4
4Vbo0tWmxS9c5XvX8pzssB4BePAkPBVdZXs+GuSjXRi1vL1D1YDjsevp5hiqnRSq0pTHfXlPwmMj
2wEGhXf+xdIaNUKtgNYLAxhcbKQeJcqI3u4WgaHXeCj9J+CnZD+wJ/vwq+s+WHCFcvuOO2V0GVZg
BUKzcxPTzeUZztAV7HU2Orf/3mHKODOY6q8LlwQIV+zBcpYUlErmBIQUFuv67IEm5tKK96DQSYBa
p0nL5rHU8/j/j0BHouhzqc7/pumRUQ1G2ezA1aYPlR7SshUxGMp9RD0FjcyR3XKBTbBmDo+xzF+k
nU1vi9Vff6HeKobYhFocGPhtQumP5GIRWFFda/steT5IkekLw53J/76d+oQDGD2tufw68skab6t8
s+R8x9VJodVCIhDSxbw1buCFQyoijuboPkSzpauO+w44mTAjFQRQf6bxTK3+zQSBfq4RAq0RIxiH
rWXCryuPFqKDwyfvRp4PPGNxKqSlaYAyM47PHWCVLNwV/sRa8+TiRGeVL3a3NMFMESx2ryZm3U0O
rKTycMJMWeZy3DJqduMjcK9J+v6nNrYz/2IbeyQSw7IgRwp5T3WeKkxWIyH/E4Vt8FSUg8HGtd6F
JeEt2uPIx1tlIVdadwhh25pK2I3GAHTbXn3KHoo5aX2fg2gyFiubR2Sx2w6jbHe8JKN6IYBjt8xg
iath+UMO3abMo+dILQScOTMQUCufZ8FzCZL2w2UCXYhrc0IHABE6w52hRKlNBeniOalSy27j4epC
DpoR8JitNJMBZUnYeieUimqWqW1LeeSlnoQyfr+E2+Ivp1kzUx2NV6y+J+YMXiNeaj6rfy5RKVNT
NKKhv4zKoc2dPNgFZGxeD+7Ik/R+cURdRLQMsB9h3W0Z/Dwptst1Piu6XkEoB3S7LHAHRsw1z/UR
XEHg1LdeKlPE9C2gZnLMw39ScJneTYuq1hPApXtgkQqZ0FrENJwcYeU8+9So0O+4ntcz4UEwNl2j
+y1Oui9KLvWzX+Z/TrW+8LAdAgJJWhgsNYg5slRI6GrHxQPqF9jZbSuhYHPcbd8IdrOLXUcVvFDW
GMFoWBz0NtIGuAPAPUJ0QT4RPZ1pdtU068fGNSvr92J/wAEgrUW7tw3fwbAJwA0gGuB16G1xUTBF
f/66guEJZEZpMfVk6CUjpeTcw/rnGEzANNO+DRbViOr2CmJGKu8OWeplT5u4NP9cU1I1LzBjz8/i
8fWX89MFradvoxDBi+VHr4ofXjRdWg1nd/tjDdHF0NOkkll8xRKxg9Gxces5SFcVKR/HOlBIyeHG
illLalavVWPEFbwVzauR7mlbxY5CKCkztXQH040RZuegCCW6QUvEn+yYyLDiYsNmeM3eYjLRpa4X
p744y94DztJonjwJb+sW9wTU3VZKqE7jG5WeHMQQ8L8VY71NDFsi15x/OawxPDmvcTjSmwe5yMk6
Sc8+XoNb33dIHnPkIQTCr1BZMbNXsN1/w65Y+rYp3AtNyYeKnwL5Kuvwr10iZurpmnhDrDOUslWc
yjtldTHrumx+iGoKnrrq3mEmaD8jBy/9VCqqqg1QmMONOf1bUVB1JPw6tYQIUcpaEjcpDZa/L0S5
stteXuSbdOnzO3GVFX2olRIxM5FnMpdwVZqbBbqejYm2AUyP69sl6OLbHB2HHcHom2SRBDMHMiKX
vjXt3BUAAd6QVtCrE40jzWQPYbWoGGtCXZ5Yz0n3VVb0qSUZnWjVfmxLC1VbsVcg0wsxQ64Ko1R5
MawW8oKoEJbCUeB+YKtw3H7mrpty6hFvA0P6I29pewP+7xrIR6DTDhx56wNG4VVQsSLRe3aqgzcR
E8bbA3Z2cjiIM133pZWPBGwa92F3S6A7Bt/WUr9VEs1rWNpXnUEhzPoI+iWFMWCbg8OCcsrjIiiY
gShWOVrbKDF8l3Su92JGntC/bxcG/vfPZmiTnpgA3dPhfwaczsocMivq5TWzBuXKosAxflvdMwRB
QRyzT7y3NHE0Nk9j++zLCEbsmjZAHllXlOjvYhx6eU3SiQPBs8IculSsHgidDBrEXOSURR2iDpQp
JJ/Hu9gQAvSDe+FFdme3y3Lb3WdtNg97Jqt2TqWkuzGVoDYrAXEjJreJiPmgaKB2Bz0zmW80eBEc
XoSuRfNEzFLovsB5TWGyp0icyw+EAB/2dZSUopChK4PMEsjVQK59YUgYs58Cjk6iQLAzcic7DwYk
g9yVfFG35hSb+9suB+8T1pqYFu+DmFzo+tCiIXaKx8GsXtgH7z1Xybqj/i/3aYR2gHiHs2kQpQF3
ACZ49/yiOdjEUsfdCklihsIR3nZs6LzCAzvgrNIwPIVBKlqyMoxwr3S4zFI/Y3nhPJ+a6MOII030
6TvsjFoFGWMjld6B3B+uVC/btZ/VSIAyiqxMj9UwJzFtqonjeEuzyOWeKWllaCHMtGwoRpKjWsOV
kZD0cemRbw68ZLePVEd7ijmzHRdGQ/dGDxXWVo7b50/Yp/7z/uOMk9tVBsglgo2MjOt2GrUrVvFO
JMiaWsN0svcOPSQk6SPhTTEh5SlUmGBRiz4KFPiae5/wBArjf7+VA+5FFn1Fy1LULXtVPm8gXBuC
0GV/XuGs9GDpVJ5+n5eW5wxb6eRGNvrSKKakkb2qSz8/RPoKdIOqIrymZiEt+IeVXbpN8DVlUGnr
rb/yq5BxCBt+xAhLmm4HS7eUCJlPZY8vRZbQswWAz90rGAZ94OoYbFMVxkPPvok10066IfftuNIj
lzbLNAyFgZrFZq07t8yoO+kIae0RsKepQGlXo8Vw7LtqymbkzkTjfWjywJlbBE2FhHv0qUVcocIf
jzPr2FIJqtlbb0f7qi5btbcceLt4uDDggzgRL29gGqDxtWf4CtrY3pCA5CuyLroc11krxzF3kgs5
qmJfLb3xxFD4Ocq8dvw+r5ctaC2EGh9+fPgcZ4YXejzvlOsibAL7py0o1HrkfPq94Mc806eKQ6ch
tEkfRd4lbCfVsddVxLA3dxkWaigWFnYdzk67lMVbHmGX9ipsN26eS6JzZlPrS7f6BaVbt/n5c2tq
tVRxSt6tl2WYqMb2r1CQLey2aFWDqCeQII8FjFeJnXJBr7FGPxysSpe7IVKMXarPvxQYeIGgfQXF
6BCiE6NT3aMq5cp4zmr/DAipZvcCv4yP04Ft9eLGCxUyrGjJNXlSvp4iFQQXPVVyN6P9RJNW7d0D
ZgoYShA0bEc/Fw4mqqkBeC26OVY1u7noI/YuXhPxEqpVA99bvmaB0q+SIMhi0OpVMx7NFPI36FUP
3UUmaOLawAeCU4wPG7SeNOR7PRR+AseRV3TJ0kf/4oc0tJCBJSHEu7igJFmX336UiBs4m1OA7ien
AnEo7N3Y3Q+h5k1WY4zgUN0y+x/Zk6GdRuLkNf4NYqe6dNd5q/JoboMNuqFoMyXI+0cYlSJ4P5UG
JheJcsPthq0Sgv3+8ZsOVTvKsA+C87yjOK+P1Y2Ww5Yi0OxSXYnSnIHPgroddb0sntn15rVM6daI
kzEi6YhQ5h3ihMDY5/fESeCCho1LckajEx83LKG0te+rWIT3KvKXlScMDZOE0gPxbz8wcAR9Rh55
We+IRT4FPE+AIMEn7dLFUNc4tZPMcAMmqNehphqpPjyu+tyY5X7aMm0qagWBNUrg8+/Wx1nxgPN+
6b0/FmARDXB1iUXPTPPaABUUjflfGIINjyqtHoZP7ORc44FRT/U5Pzm5RJ1v0wVR3MZSD7qpPrfi
8gUGWCwvxlU/TwjOhlycc4PUALYIulOtOxhnEq+UMmO1B79OOfMgtZ/t4L8RqClouzCbLTHHpT6w
YZMt2cCzcY3kvCZIVtXgx4cXw/P0fkKx83szoxFsL1VY0HUElr1+sUc/ikDVE6j3SohYZ7Pwhede
QvQwZ1myXAjzceYGtC1EabZSOIiP8AypBng6knBEkKMxr+CniFIvNM+Zbst7bdWqmQsSZVKTvfEG
ruVrjHkbg/Wicjw/akGL+45KFcLqjhFfs8OcCYJt8ES/veScRmBeU5lihu7ODUybioGlDtkOPgBo
s94p+pPoZGfLPIyRROVvuBjA+vhJiDxvDF9hUuK53WNO7Af+DRf6AyXGkuHTZDYTn3Pb6+e2QvRF
leKgGffbfRARzQ81qtScWj4BimIv4bYu0CNg3wk/ChbwFoZxchwl7azqf6nRYfyO6XCezA9by6Bj
dXUEPHWoikCmk6MIrJxoDgOpnAOJb+mW4sbWyxaOukDJeVQlxY625HfiZI7pMgTuqJpblO6l1YuP
NCv+gZRoR+A2XRqyqaZIrbfapuNlNMxHIPOjw1fx9eusKavV6CMZ9r2dyZPunnvE6Gt8pNlQy6TG
Ti6xZnJqr6jGktwr/r3pL2gxUYQjFgowbAxuXv0AsneNg6uQrWsrZlr90H0TMA9RflZzMmcc8gOZ
gD5X/4z80bz8cm8ooUN3BOu5obCoRDyXrRUxrqrx8M/R2Rje5frA9+YUiyq5ZTTy8u+8lTQv9XOi
/nvwJWsIMX6sauARWFqIl5Bbi0xFKQ7FGS0Jl77L7QxuDHQ3Sc7VoR4DEw7d3SaSHJ1Qq3LoVyKC
bJfHM0vvcogtfeSQpFtorFpmTwp5qQi9E/dBs3IJQZHx18+LEFiyAzE7CxxyjXi9/JS90Kc+Fy3q
CIq89PMy6VvTLC1bGErcyjD1oC7AC0iDAKADRHezKQY3xSCChNr38ysRoBhs7Hs5XcFu33pYbbqe
Vb7FFeXLzBRKo8FE1RCScXa71YG9mYnmhH4gp45m6hPD4QN9QePgtXrq0yXQcoQTHe1fM/KVggkh
BNNxu+RXr5UpXakfGPIEoF2GM4AnOhfTOy1LnNDK5Cjt3nLiU8hdaWf276gyfXEIqtGM0/Q9f8r4
Zia9F8ag9CL/nPBtfTazqhxpeeWxvvBMtV73ueWRI/KAVhYwUcm6t3EuF43Uo2AsTu8yTefVojFu
hFe6Vz4N1KVlJEmz6+1tLsh9CCwVgEaFr8Im73KfzBndY5oLs+oQx2mFQjgfVLRSqrJnSKWKrNrf
X2fcsER4diFZfoDegWdmQg8K0tHpiSBRYir6lrVuf6oJBFq7ikwu5kSn9SHspZm1EZ8xcVZjAJGS
nHeDmBp4pq5Ir34e1ys84v1KvrqUM/oFZUKhqPZvE85TZoxtT6UNdvD/r451UbUw/3pM3SomuCXi
50Zw2Xw9bSBxOtS3fMalCMv+pqCYhUzpGZFcIetLdkrS1MsJAewbNCa9ynqvaA5C5W5VD7RyIfpc
ptvHAM8/PJjAlplfhsxAS21LDZxRPoDX2RYt0UicZLMQrTDkI1ZwpEYZFNA4UHi7lRnFwATCTNdZ
2qkXZw37bVSrWtSwkWofAZcJ88HCmrUBKNQMHiReA0aB1voTtmLZD0DOBcU0Wjx992M6js4sxC/5
pS8rs+pOgt4BzhQljmxClAfgfhFuUD+sia+TwOiNIMXx+gTO8A+uDzMmLNpM5fTlZrhkDX083tip
CquTToobVcLF3MC7cXTdoIIJvPVRXw0mWq4sK4ced+wb3WbM6Z4DqAah7hNoj9mV8JqR210EyL7+
PcK24B5b9b7js6grLuQ7WVsqd1UZqDbpI0DNURVBTVvzAZZbxWmo0QHpcOUJMvZHjYvUQBugZk1u
0TaXa1I4q2cypl8Xrk4ueBkKkTMb3QvyXl4f5SVijmYVIg58gXkOSjbvoXD8Ie9ugs26zqvwpPch
E0/nPNzyHbCqKjD4xEaQ+/xlEtmHF8w9mFpFvsWH95M4qWUWa21YLIkR7gJdX8y3L/Tp5KIZwLuR
VIzyWawEtJerR42SymdhtSA/I4oEBR0P18PpwWGxZYUXYOgtc/OQIVj14E4xAsv4VzJB3CoRjwvV
elQLKPAnu2OqDLvP/b5gVejhwn4Un5Lb30ReCtCgEhJnV3FBDCpxzap2lZqucAOHfFwQ5h36pCY5
fdox7bQ/c4dGZVAt7c7mlS3UYktxngCtHH/sxxbGSvyl1hv+jGwcAhNv4mUuruevj2AJMKLvJgU5
wXi3nzkvRknyTZU6s6Gs2AQekxyrXL66bHWfhIsCvlB3cL0/80nXolI0IVvPKJddkAzCSajqEbs8
zRHx2hwfiySfuWuDiRo+7rqSIWCGz3ux+EyMGNMN/nG4Rj+DLvxrSrKftnzRkL+OnvvVU/sd0umV
jG7Lgs3cfhBm1MQOwvnNHt9OTNKegzIIuVltqSOoQVvaBNwEnHJvUsjLRBwHBu6Ev5FvkGOe37IS
o15fOgUXlvA3aMiDbxPBNhhKVWH+x1rsmX6+GglpIKxLN23BBFc/2vrbw9vXr3jUILCHbGakBPfD
QKd1FHXkPgNgaazUhzyv4DghsWKmJ16zth5Xe3psZzeZs7QAiqeDTyXjB75KDR6lWxMVLGVWn99M
A9ZalOKYPFSj1e2Ri1CXubS/jUR/XWw3hMzAb1hPEOi2vvW9mEaih10GVcMx1dcc6LOqlMf51g4s
IUFR5brHiEx8dSfFznr4u2W8VourWSqID4Q5VGeU6XGnUUiAuCIeu+ydBCtYo3WWo2jWluSwlD+R
73KUbr5QJfKASuJEO1iua6v2xKXqDH2QT92Oz0FbSWlVwRSgPYiD0PCDNR7DJZUrfTHaQr8V+zEy
6n68PVe6GsO+KOHphrnD/yG3hOfC2RJLZ8vw2EGwxLYHUw383slKFIT99/z2YUOXNuNNzcPJKDLz
TVrFVbVi9c8yTtG3rqg7Gm1Ed41bNGWOE0CrMOE95TesLAAfWUwqDtahCQGI6RMtKbZcVjWXEyMz
sJWdp0yqVGj5N2OR9Q6yUsk9SjYh0qmyIukVcEvAvhQPiW+tiNh6l+ynXe2Z+DJOHMjmBam+9XaB
lTjgEb53XnKGBV1mbQCMT1Ihgboqmyq8047cVE283ek93qIKLXs2sPXLxA4OIQlhLU0zU3gBRq05
bvjNZItORepIHYGRVPLPGp/g8Tf8We9yz3al9ykDqRpZxiRiW/tykBRD3PqWkGeCZfdpwcJIInLE
R57waEIX8Jold9xbb+Yxod3NFcDxUGV5W17P/J0RZWQ6+QSpR6tfr0dPgynmZIV34qPj6aotoZtZ
gxmaAIhs+DpoL4S2wLA+4QpCdSYISLJh2oupRU6xRLKjtPNAq6acPO3a3f2sDMFenPVgLCY54hBX
q9lrHwiDp+JQ0kqPqETZqRmkspKmIYq1dXHkFeCQ/ucla1lQtC5pt2NLkZgA07hbrgA6UN6714S/
fggnpgdptVF27wEa8llKX+WaBwgr/hZnMhPevubnFXtvMSifB1S1e5VpBNjhgFAGlHNY5lpM6VJ7
n0+38idh/cXUvELLLThNkoAB9DH7HfnTqQxSKm8HQds5BNQo9JX/1HJG1joIg+3B/x3ZRlhamfuf
vCJwxGN5WZpdYvLPM637iGj96e8BLiAGXhn26wpWzEYGFzOJjy3rQob35WYY+EkJcevvk6R5J80T
A/SPiiL/G0XqB5MvfXkrO7uROW6TW1JLCsbWenGKbzNatKrAAtnCXAdj7Rm3jsPVbnKhF9+SF9Q1
5YDUfQeFXJW12aHlha/qFdOvL7T/v1o7sKdafx97U2exDT9m0eyN2cwtsfZOZbBFRvzuDLAkFl5s
IV64Iis2RWQqVu97wpVPpcow+38j1XVPOmjMU64UPtF+PZy/vYxdzwLFifiWeBXnj9WYfsPEN/fp
N1hJxk/wTpL21KslCPTr4pQPtjYBRoTh+T8irDnHTtg209U7Pe00Yc/XxooKMXgBP0ZYn++LOT+w
PIWFazpn8yNzw1QGVR4zxtqMa8mRlNBokuk0pvi3TNr7dLthkFvWkwtPgkQrOdeONF4Qt+FM7wUC
QHPkjfZkrKdoo1GSZBA7MPJJbGLt8jm3mcez6XRUUrtOIj4rAaIw5ydmplqztpwg0fkHCFeH9hz3
bQLkd8PnV4Zr6fN2hRRCy4cAS+cQoLGgc4KXd6TOzKvmsmBvs7Tz9YXHA2pN1uw17e+MG2kLzOeY
gDPIzCWua8NWa5WMti6mZOsQLmNqPrkKUPf5n6ElY4sC8xRd+E4w6+pPQpHKgRvTMw0r2SFLxo/m
HhAgro7sbWTEwqjuVwADZcxuc3ovVJPVroSXCl7qcIci0bF1NPqCuKjPaaql7ZJlLkuVX4IPpsvl
OkfbrHDEwbG9FUh66vMmbMLdDutrn5Qqhmd2bMa4F2ULhlnNOiK4a5HIdEFzVUOLr3h1YCYH3DGl
hH0zg/BpTiABO6KYmVlvFPpA0eZawGT3S5qQ6Zd8cgC4Bcq8siIDO89bei3JuInZkzZ/mVxV5yo5
pj7kiTESLV4fIEjIZ+u4G23Dzb+vDdF/eCVIDiWaZOMzg83BKD817J2uHKpXumQ58578zQP/Gn9d
t/TeVFZ9BFRC/2MyT/o8zWuji2c9AOG1fb/AB3Q0UKKHBX1/eQza2LGphAVyPT4woZAKRxpn7xWT
T/3bBcfvK2QE69+1AdETHTOX5elE2xsiaEgDFpyvxEzJKXuckLp+FiEbB/cC3XQCT56ZmCe5OI1A
rAAYKcOl75lT8xVRXykMvAsz/YnqBzAKAlyNMRg8emklAxe2zqNoZtMqHjrJOuZYTN4+X5Pbc0Gl
w8NX2wzmATI7y7/RDIIDI+q6KmNlLGOkF6Ude4/2q1HvFZZ3n11oaExxWMNt/SlPCfk9mKkUDgvA
Hqu/aTJeDFEZ5BQ2WibKfr/hn81xb1iuE9fFkyHDqdkpQiOH95gUj8mh3LYTR06wBXZB1U/Mcwqy
yFQg64l09cenXlsQT4nZ77E7xS4sQ/oOSKBwiyIzCsLUFrqMBPjYg+lTam8OVtrKqlGaY1HV4BZN
qbIojwW8FbcpJqvjnOC2A9jYE2A59b/27GudQ3Z+WLnYXDPRxzVeZyzq6aIi6L+/zHe32e/Ih/f2
Jp7MKzYxkbiH1h524wuRuK/veRDgLNiYnSZr925inKaI0+7I19KcxD2GrduiTEy2uUMjf2ZUrqj0
J/ImLxlcXdp0oEnVUrzB+bRsYoRX8aX3cSzpiq8deqX2DXUytsZX1U92crQet5ygopjf9aCKvbKZ
6JczOCNxCeXse21BOyiQskraloH/V5vs7o0cfVIXVyfrirCPPGkeygB/4StUdfvD2f2TUG9/jvux
S7jybpC89SSbPryfzL25q+q42xO1LaFuCmJ3CfgYaRHWTc4bwWceyOwgV+EK1wy3D94HfGXTIQMx
zo+sX7jZ00kc+qd6zEeAre5W07a0cnvy5tRFYXTYZjPHGxvue4+6SiNMJrOlaQisYM+JAeE1E1Vv
I97itLp/gtQWvVwk+IE+H8WkMVM5fliHBUaC2jeXw3rTwo8quqHjYFlc9Usum6zgj5YN7mj6WMsn
wwiPUi/grmTD6shFDzeGArY2vDNArC5sMGwtiXC2KhDEKKOlQEhyWib3bLFWcHXZ8N0z2mbTEKgT
NxivE4P8/A3K9bYx+tkep5PMwyWDCBka3gw2TM5h2V++xNkx5R0K6vyc5twqT7ibgHzl+9Sfw7RD
U0JC0eMrU1qUXj/pp80PpWdw6nIueOW/safjXc9Cc3Oz2yNi1xpU2Ak5CF7bEcC3MZVtTMLhWIAe
mEIXbt2PlfXeCTRFRQ4WPA4BrPHs1sr1WiY1Cvsbw4oCj0HhUKrv4Z3vGbu0vCIZzcAVxXQ+ALdu
Cxb5+UwwE8eS+n8rhftTGy2TCJIqJstsFlX2HR/Odus6uSkT3BP5V/ScaBGiBFd3dWWKcrRJ1765
IWQYZ2vUQydvukMRbMA777gF2A2VwuAWFyev4aj0IUBXtzDnuU7mRaPLoYfOyYFbtUokAZ8sXP/w
o2TJ9F04QHoanLaB8h2f2PB2FCvVWm+/78iRRjxmgEpJWszMleWoFGOeeFDYuHZO3c4htZNv4YUu
tpyCpG7lDcwKhtzcmXdH0lKogODlk2+1h5f5ijAWQltuaWjEVZJjNJIy5XH+D5jCJxIRtwLRnmw1
AfTPVYeoHuNmc2QHfB/u6Z6ReSfiX/nqxw/RBFaoEIbficgkRlwziEuGKRvW4tBdLazETeE35pZs
6GilOZKwiXAPJt64kPhJrGtOKT5D3CBkRyfNRBJavTfs1t4xkz8ZHxDuuSMQaukw6e5E8sKpyi6T
7qp73NIshGZOiacbA+6d8azgJyZRZb0jhO/Hx34nnihKLUwd7BoROUExJpZ1gVSKWIxaM8m//fam
lbmhxcmCJ0AWEgWl/g9e7iSP6eP2Q4rCckAXyPLu1xVy2bIn9bRIEov7AsW7UtazBkrQcAbDhIsF
jH7/lDN4RdWR0NGRgqVJl6pFtmR3ELAbI2B4hJu8bt/aFxwLf3ZcOlHVcqS90GJN+g9BJmR91t2m
9HBPiF8pm1q0NOoFw/RmLx0H2fKi3yrhNc+gDcu/qQp6R8F9MWuyBlt+1BqRgmOet21CwBAxyofc
MulpW05v4M00BLtL6tgr66NNKQJyAJB/vpc2ILLjuwyVvr9WtF8NOnhVQT4EhvK4zX0BvUGyQADh
MxXPYmfNqAtrQ6jTKV+76fjIwtMkkTj+cXyKI+MJQYi8KxXTq9PM4+S0o/qcqDrW91c7axtKs15o
iZsloaSBGhV+aBsIJwiIq7vLi0tcATlDCvqjN+JTyn2XBUGz5NRv/rihp88b8BtyU3KagAvE1/LF
h5Wg9uIOwmIWFPnnWf2F7e6LUouapBh8A64SQnAzMk2EBEsV9Wgx52nBNZksdsWeioU6T0syvf1c
yG3HixQjIaxUlVat75QpV7AUrr3uxn+ZmjxV7Qx3KVELgwkVAKiTWZeD+CDaywtkKBqkOu7SQPIH
5Lo58gV3op+909DYSl6sIg1QuJkm6F+KkmLZtmmMaenTLawbvTWbicHge/5sw1+IkTRfLMOy1Q5j
6Aw8zl0tJZADLofpR1Mu6/I63CVk892ONa1fjwL9aep0iZOmS8Y7M8r9Roj8BdRvseDQhRqRGU6f
qZPuQSm7LnjmrYl/ATztdFTvgd67vUqH1TuxFzrJoRvLZncwQ+XVn126KhZ+YZ0JFT1hVHd37cYH
j+hJia16KlcMUVPFA6AEdXYHtMOjXzQAXGYhHNIZEd0gOeR3bU11sMrEkpyFLdgnS4orbCzSjbrx
UL8HdOInLP9uT8zBF98PG/k7TpoXE/soWiAmpV0ZxU4ecwWZmT63OkZn3HyQxeX8x2Vzs+wHJsN8
kyWp4Paa/Ry1PtOAPmMDMjlMOcVO/Ke8hKVsviBQLim0T8lNQ1fB6PxSTzJpmpFNgiTnNi93HFtA
SH6moSVCSu/rCqX/AWOR6Ti47G5vd7PT1CU5dH2wDdo5PMAPZs0m1UTtP05VSM2K/q2vElqDJcox
pZRfU/Q66hnREBHh91lFVQ3xOVODXTOT8xWGBzlEYZtxvNw1L/l85h+iPJckmMUkPdihyV/yqWYk
3vhPpgLzScV6VP7wbvWOapGUzcXCpItLY+gtgYhTyuLiT2Iyjs3Y4E9IvOH9qO/Je7DXQ7ABfYAM
7u8pej/K9L2twoCcKULBdORtHG62v246LCPdCYJjDMUZ3BgtIjW1JZox8ZOYskeoBLeL01SQzIZF
BgeE3ue1C9BqhKRyksvyYKwKyxmVgnStID9PeKeW60C71c5Ed4NpOCdC6MHev2L2fNGBxfifwxsI
Lpzz3GcLgFFEjefLv8Y0oSl2iHvEKh0EbF8mo6fISN233bOluXwCI3INNXvo5ZSAgPX2I3naIKbu
FoF56xFNNwgNLJotkijrgXwyJMtA89bYOzK7MsIpaNadONCDD+Oc4mIQHzqSxStmli84E4CVOTSy
/wWvtALzRo52d3pYAzK3TALhbLSFaBf2h6a/ECL/Qpyt0fiKmEiM3M/qB71ASJhaz57fVY4I3ing
2zoQWfsVzsXurp5u9YP+2cPoqWPnrTU3dbE66YBalSQxggU+UutJQ6rw7qpg/5cfWSZZGiCqSquA
ETEW6WrCg9uTxB+Ak97B47+76fplwsHlZgFtb/lqJLpmhhHLucmPggxJHHt76WhJ1PSLe3CBL2ZT
Eyaa1X2JSngOk6Z5Q+cTZBPxIo04TFDD76g+51yl9OvG+98YROqt5K1JVeKYgez6iSwtJkIceN3Y
0kCjZ6NmGsVn/mXvXX8iVMX918+mnnldE0os2MDr2vwznuXYCF6+jhudETw/vGivelTifBNNyz2d
NvxEjTfjrJXAVWCrW3zxoUQi9/V4naDqT4vBr59oj9j4Bfq00V4fWLMgRiHlIQrQRll6bGbvT//o
8KoGnv3NwPD1L/pt6nkOUncXZPShwBAuWOf6mUqRBKWDDHMiOJ5SSoaH2z8bgH/d4JWHliVaXOym
q/A4ijHDLkHE3yAF7ybG1etcedzl0tTJvZnBRRPq40tDgvMXMCCX5uaQRA/3AruisLNxbIwaxEbb
DiDViAADG/STD7wIJFLI0iSJB9iUrmS53aqX3jBJBFAgPnYPkZ0cURYQCVficrlhdFRniadIOAAD
WMuJnyAFoQzMJfX4Lp8YzoWkphfd6Wjo1DgpOipRRO1o9DtKr2uy1Zcaxjz5ChhFfiWKyA8hol7K
I4yrx+gncM6BpQ9dXlLYqe5yW+9Sbhafrdw98btg0/EppuqfHc8r6iXvJIqqeXOcsFa2awKsg14n
O9AnyahTjs72YKcslyrkmBjGlZCATEVh8zz0bU8mk1YROG0+rsonHpW1IRelEkzIc3BbH/jHGorl
L5I59bpyML6NmcesbcjoqPXFPRD50MtHXG2zw2RQu+Oh26GWjDhRpxJ+G/9DvFf4TCwA7C8Fyv26
9NcyfJtHLobGV6zSuZzgRl2DaGExejs72ZB4LZ/Ar3oGxVzhkWEkAzJbkf8lNd7j5v3FcvN/2iri
ly2nUoGs+sMQ+GQ71DuLRo/D04NYb00CFRP5YpxBZO4ShW6M3/XSzoFJzfYSObUpc7vMEoO9XGxc
xgQEl6Q/rScTHEOL5mu763oap1NacclA2jRKhkP74nDdaWjaS1yx5XuDDMWW5KTCF0iWewoknjaq
UMwb3UIl0ag+wxxs8AgyoXCzSMl4s0TKbo926ixAyLWfu9Vd4GP7/q198mq+d0uiwl2lVW6+WyHK
zh2G4Hqs/2hltXuD3vohx2GgPqKloafKAPcE1QN/J+nGBAXIGikjAXQJUvjOEsVZUf0yi8iReswF
UA7uk69h6bumfgayEt4qbd8DApziyt6trPmY48N+IJ7sr/mtSJeH/1vTa75zSuQWrdbagfGHoHYn
g1ggOgZmdmcbsynjfjk53YxHEnbJR6qw+K6y6Km8FWGCAzbdgdmBq0WAN5x9W8DNOt7+j1SGs2yx
bzzNGTBtlLZ+ujDQXbzhnNwrjYjIxPSw90CsBqTI6Oo7EB5IjEQj61eRL6+vbiWzAIO/GKzdfr7r
5zAzUvTQo7upcs1SrH1or4/Af/d7YXTksaN+ZPN9ZnRT3qGKzNvwJa0nIcgk8D/KBp0GbIXPeHri
Id4n5twQzKsgDw/zCegZ6SVecVq6QmukZsQdz90uXJCqtP8CpyVRz5u+mUx1X8qkkID0cExfIedv
432+0FfNRFHQ+tBiUHVfiwbqeMfyZGJXHpQfpAAX/15n4bjofJHiJOcuhviAaMtSZ305aMMfLpGR
O9/Qvh60ZQpTkhczN7iOtHQYupKuPCoTd7SLMMqC5oZJqsV0utv/fVvWcyFd4Nw+N/7aqsKTjJSQ
gSSrJI22AzyYv/C3f1srrYDFIrSN5TGzUEwNogwth0UOePFYGF2P23MJedx5eXtLXj6Joz97pSky
qvdUlZJ632BGzgiiWCjrO8tSrDGtxDrlUafiIGkq9ZESjGnUvlhUemzYMGD4zs4+QJiPaI+bJDr9
jce0y7P+gzAWzx4WJ1YZkEpPbjjUoNlR4QxDe1beSoOMX4qY+0D4UetgxYKYwEABMe18dZQejozw
ZM541A2m87ao3Fiy+F/0610GoPbfjPZXQi9IefMKT3GZRmntqSboQtzqu5mB0JjNHufbuX9jlIkR
7QEqcoJvvyzTpx1pYYFLrw1jH/JZM6xgmgmaB3qtqGoGP64FFVHrNgeHkqFgfxsdZ/tDYlmiVMMy
FLpY//js0goPNs1Zpym4ESp+0YPAOsq9HEZMOYG1br+zHbj7bxhbf6QKklfGb4dnEGpkWtBjEVEc
HxS5EP/ARR7mgKtY0fUTDZzj09ZC2f42sWiLrrpmtrUtvii9jVPAGJtHuEgI4CRf+tqfsNiiNTTI
YqimEUgjiml7IH5R9hMcSik61dYGtk7xJp7QB5LKcWcvThxKQvXSV+4jyXcpKgiTZO2EF5et/N/O
1bl8eTMtLxZSDmwbove4ZpwF3Lf8Sv4d53JOAdAkMQd5smYIbNQn1jnNNtcvWtdTt5/7i16Arc0U
XpcZUpNArDcFYnOM7trb1my2Tr8+XE+/h28SVc+hdeuNASk6x9pu2D4nrnMt6oAIzSZv+pF/LEQ3
E1XGOLo4HvnMDsahVZxcQJLQkYX+jY3XV09cxRSUoYpOWfzxGOhiXs3MkLL/ad3eG14Y/D60QRKh
k1NVCcwJDhYiq405xTXgyQAqoRKf5cBVL7iJqKHCSPvIggDL5Q5rxyjgdGlTgG6a2wFsjXKDmhp6
BaoyrSGj9QrdB49TWird0Zb1y8usxOxN5+ZSRF1lRVieTErhu4akPQinw2tPd0KGImHUJDjs4sOF
0bWgNwwJY65OU00tX8I3ifJ4V4N/MRbyNQRcBcBUkI/KHhVrZg7r3jJlLq81MgYFWQ/OLuamKzjM
gMWmFO7P+0Rch5Hclkh2PZ8kTgdnc8GFowIL0z/kn1pzUGV0WBYkmqED5KKHbQIMhobbG7q4mYGB
39NARTXaU1xt57VAJOTCmi8LmgnYziUTWpVPh9fa1ZWsJdAykS9A5MkSnb93dOrPsaW7WFYzgeJE
VZXsTi6ZGrrUcd0+G0ESH2EooSWm8o4NNLwDC9SswCjLCiBhPgl+Wf3zWlRxalg9X8Ao/RpzbCxp
fFJG348FoDL+hEVSQjFv84DXvFYBNvxCCtCK6U6/DtLVKfXJMoPFeaV7l8qucCqeaX92UkBskEeO
X1RcUtzz8rjerJx18dPZr2jie201PwASMFq5hNOaUVJGlClEs7w/2F8FwyA4uKCA1hOfPKLbFaeD
W+ZxgYPMr5+VMBy5Qm59mZvkJP3lCSX7wbGBSTIw9hOV8LIXsfpLoLfCvwOx0v0WbPAvKf7XrBTQ
vv9nc6jU1CG7mtYxbMweX+YUu16qWFF1ob1kAx7O8aNQLo8992Q4u1n15NKEbaBGipFdx7TQ+fe7
SYV43eNbPhpx2otAPkf4RVZAtJqYQmkr7BBZTTGzNGw3Nlu+9iUstrpxQYo8tjlW5mtTH/nBz8xo
R8bb0+XtrUAFq8+zEBUpxgtNpG1qcXjxcZgkQeQH9x8a+UDruDCVgxC7vMP81p9OnEs4HO5nxPwZ
gsyICqnrX7sODqu1546O7BKP3UCsMo1F+XGhUG12A2irkfTOUfSnMgsZsaiMJVRcqBAqHo3WK36A
clRhMV9h/n2L5RKVwNBG1ZBe/S8uDmfBB+IM/u7Nw6YLBdJDcJzzsEczBiWZI/l0iZ8yU1Zi+75G
3a1iH/2fz7e9y26J77zTQUMR+ivYd3CO0H+rQ/7ikktQpoklEIcVX1NZ5mmdZ1gOto0igEOiY6wg
vMcy+Obhyvr3EHKThi1ptVjf0wkdU5DijfyLFEH01I+3bO31KiVuaZ/BFFkT8QiG5btXW5q/XAYH
Qu+OMCLFy6QA/RB6gtyt6hzq6dzK7BGaHSP/uhJDeDOXoMdazH3K2E/l35XjRZz3aA5eMaUAJOOJ
cPycpBUi0WmXpaVXvaN8SwIb4NergPyX4WKtOS2TI6UenPMRdLwaF9etMRtxKO6/zvstjlCBgdeA
AiU1t00HrAghDpG39WftTBUWT63euJjUH4bfCu4eefSwO8EzFopqCc5K0ZC1QY4EsfGqepafdQNO
t6q5XsCVUuolJnFkwm9SJ7/XYurJWeDjivQpWlwflVUm2V6OYLcNWmVaV1elZSTferlqRB76hAxU
FA12m371gBcqN3RKap/C9SJb2Ruiom5zaCBGdBG0Oe113OdSZAnO1S4/i5ya1I9Fl9AMGRHJKvSt
4yOFlo9oy6PKz38f3QCpWKHmN6ddpaLZ4im9pHIUq33R22kP9YxzAxaxXI3Hnm3Th7aqgMGFeNVy
5Tv2mtyn1/zQ+6lK96Do9V2LontvZuHTHBlzXLhd2NvOY0LZQDFvpF5s9q8VkRguC+J/OzsRycsI
wWTYjnpY41gNVGjacu8EPvZndyxi4jF6YEJcm/MYKQpnWH9xBDdwxP55u4Vn6Pyb1Rpd/5sLRgQP
oTp9J8al9JHY1wQH0MGW+eGtfpPII3A3M8/YtoTRngpjt3r2QIAFlBObnTh/RY5wuRXUQpO8WJf7
o/wHmPRkG8e7ITVa7C+MA4t/ro0IAeSxPZqe6wNhsw3NFip/KdqoW8Q3+KKbRCyyTsqZ7LLRXH+F
+b1HxgvAwqjlFkTDtkS/rGKSDzwaHZQMQp0Df/bEnLeELHBYHeiuJOp7qAYa1J5HIeWoodjXutin
3okh4vRQ4+tNg6pYL9uzJdoGmd+JIB18nxL+pxnyqqK/wpOjFHB7QNXrYQusRGo+LHOrUsvRkcfk
Zet6mmHXVuAL5FYluj29DmhOSK9ZxIOnZwVpW8O6wO3LMU4upvL+/5ZhE0a4LEtpFvDyXhKGZ3Xm
L2KnGxI0tl6Rqqe53gMl7Ad6S213ZjYwqKyennLdx/ad03A8ozaU6XWqvKAoEzFku+aLnRNqcSVd
HQ7vGtpn9RI+5KC0vdb/tUYgN63nVqvGP76UfL6zNpeX821yOea/1Rn6z+nqAsUTTiAv+OXWuOX5
hikPPpUGTbGiEryu6VPQow7Bdo9NGebeZPacOSvZBIaMmwtU3OPzPZk/u/+AWmjP1VkOt01xOYCK
IQw5IA0Dkfc0+FnAuse4qramaZDfekYz1EnO/Dh+WkcyXWw9DiLJ4mlBwNSI9hadqrjx12ZSKGtd
E80I0+lIcEJMYvcx6sFZWpUBImrVh1oc0MOlbZax3X9TkTQ22f+HVNvVgqT854uktZNKaXBW9YVS
qEvaUcH9iyo9cdxCPpBwsCinP5tR6q+DGFjnwfZrFOs4/IZUK30wTc59JUtnTC42fCuRgYTlYjEW
Aq9OwfQCLM48kmSr3Aigv4EGWqoigiOZlMOI9EldJtXdDuDdBQaScdGF0VL1eeN/MtcQW6jZtioJ
Uz6g5JSpR1eBRJwNZ1PKVgxu3QhHsdBCXazCB841hoNGWjp+2+u4/0KpdgPDlRxyhAyYHuc53Zcm
mm0CZe+eaMohm1yAGEs3JPCdWpqpApVhsqUyKCBs2w0NPi28xEr7sZtYGTVFnl37MWsH4hOOHmLc
ozkjGDmIEnMaLEsyZQC1HBDyBwhJ1ugcLulckz6gicxdsJmUPI9HtGJE+/4BfnAh00GZKtSoYBWx
4gSaSOU1gbi33jGesL8+/CPKrjgCQYEglD3cCfA8w85Zt2Mf5HoPFLyJN5SvkP9Ux8Byd0VIOfeq
G2lGLQ/NpiNGJ1loeYuOwDkgEjsl9kTJXidTSIb3QQK3TESkSnY5MnO4Y1xuppyt8Q1lWL7J2NFn
ZEY3imEbHZUq5iFusgbY9sgFVr1scz1NK7x26JeI8LQZv2PSgvMdkNn3SWfeC4/gbIlNxEcNDlrt
licr9nkPDl62z34vEvbnrG/dSHnWp1xQKChMFEF85wSddJRx5uNmzckx1y7OZO20w1htflBhsZDb
c3XbSVwSeKuKmzsvO4+foBKniL/sSeYNqRVl3fQW7Si+NLCRbgjpa2kzCtw/Pdu60um8bp/RbIOn
cKdq9eGgwce0rPQ43xQJhM9f2R0Iehik/rQD8aBrbaj3s/QF4aaYStbYLKY0TXOnENqeAQ92ttUl
fpPZ4HG6WLjCWkvowV1EfOqNqvPHV71r49G2pBeSQBfR4ua1xixTmD8DT4DQNTGwA//hkrGKJNgx
hQYxl0RzJm3f+d5s8hPtxrq/5VK8fYeyU++ArszOMuOvj38H9elfLuCfYptRxXkOTzahyF7PgoUJ
v979b4/qC6pas8nTKrYyzpZClcbxdTtRHTT8dtF56kfLPQDYMzcvFJMiKjV8NSxQ7jLID8N+QjEl
GpoYDebd3/g0B3bsshuGUyQHTysYGvSmE6k2/Qt+FT8uHLHedlH4GDMJVYoHG8XyV7B/0ZJAWCOY
CfxjPs149gm2pjJg5WD3yZBtO7yiKreopnjQEly45rwSASRXX6P71QTJh+Fn5iH7T2aJPAUf2kXm
ih0pkPOTnmw9Jwg8ZLRZFEQhqyNB3r5+BlVYMCb5JU0n8XaMybaVPmfRj6GIyD7wXJYDaWnUAYvb
jMEsQWQfaYl/15HtU1ZgIvcwvOLZ1xhxRbvV11narrF+EE1cvJfLXvBfGCOgxQH+x8Vf+CXj9sk7
BaEeMrKc068seZMYxEdAJc6fgP8wTAMBGEoYKIiWNUMI1VnvEvcCMB8WMTqajbYDXi6t/VKnp1kJ
8A5KBhQUh8EDLtehZF6jdkJiTt/IcRMXC4HTihlFYngLiN2AlcPjsftUXSkpvN+BsQoEUZkmR/a0
b43LP8CLhV7CNnJw1pQcfhCwkg+FF7ldNkEC9VUnM7Ap09IrEPA+mbaGlLIQgbG3ybTljbp36gk1
CwIrB8YdreptE4WK0jPpejeR9SXHdHtJBD/RIGqrFCQSZe0S5VNgnesNWG8iRRGJDM91kZtt9Ml9
bnhEHdKX0X/sRkZlLCJ2lt7vnbSuhhOPvenKHLsS+HnATDGmOjYzyaT8Q9yJ5xCDYuSy/w6YEuXH
LGT4RhoK3kKsAvenTqM8hbXvysGpwiZg/aiDzE+1DX92HN4/aBnFa9jJB6AVvdkk6VxZGDN2uZqx
llU+iXEYpoqvtFFs4X5wiOBDDM+d8yV04Yo7VEMx4w6tS/itP5fcXhl/6CzvDFl2H8o4ZDb/PJnW
NbQVoOtEWiSNj0nUspBJfq8/2bJgJhijPU8wGR0VN6WjLup/CnmQuLZs/v1pfVPIwOHXEIpqbhTS
YkO2dnWq0puphUWrV9E1SSV6xOyPZXVK8XMa81dqfbFxbTRaLbT5yh9+G3zXOEWDrwvwyGgnFixc
3jhcuAu/pZdiV1L16WNP7UhUS8Hs+TqDqXZK/Eglpp/iizXcM/eaFr8NSW5y7vGL+Z+8DZDRQTk3
DwaXskFp8X2IWM6LqRAeCYgTIQwacOnus/nTjeuBO9g+pdIHwQK02Gav+znJNFuOF7czj9r9KmxH
r7MibU+bQ4gq2Mzz8fSnDk0hmpWporiv2Euyu3olAvoUdWTbZohBKh6O/Hpd+Ajy34vDRWJjtvFR
4F2lo6FTz/oxRsGXCXVExwP803yeO21KC4siQkM0TGSB9eO3n9mWishfIB5CrjAn0WfvqT+XBgMk
eI3pNJL4b/Sp8ndeWT1fS4OPjRcgdahct0g5jgQSxy4T1OzsZhrqW4VZNNxkD5PqogW4Czj7b/IK
lYVYrBZLlDKZA3e95SVNZMGbcgLqxFFFp1pA/RLk0+YjzMk4eeMK+DQgen/UTR5flwaGOCp53P+w
awVl1XRNS60qTRgHpGKt2gylm83HCMjn5YJBy1lq39Tzll1hJeDBFtHbK7qnadeZGWWDGhxUm2iJ
Lk166wabCDir9+o1AzdXwOFaBDybTwT5fFkmyhiOXCk/ENEkoOLNN2uPIsUB+L3OZapl/bGdVAWZ
ug0fvbeTrvjlatrYxFoXjDMXUnBnaQsfzTIqTkiOP8/IyiS3nHSADRvcVaSzM6iUKnt8lyopHwDa
GTLS/XSHDBWrokP7y7a9bQKUlfJwKn2joLq6qYLgAb59NOvDUqxmxMA1uifUm9mF/NvWq8oUvjGp
buzo57KxWm9qmhwZmAWnQEDWKCNuQPUsltJ0E3JcmNOnKQSdcj/lYE2F7+++CTaXWQTCrjTdy5Jh
M4ia3y8B5atA0KFjxRToF7fkHM5qrK5L3lgzOlDx/KlKtoRj7rktLq4VYsloid62MXUa8WKsD53S
yt/ZZ4IyI0mzMC2X+3wOxSowBUlmHPXz3XSGtMqUToELV+5EgtF13P1n1K1rcLeMzcULGcWbl3TT
GHf6oop0dlhfObJwmCgb6tPIpqhs9gadImm/Vu+zSepbHuhuxgQBPpes7KSK3oB8deaknxR32Joy
7zuP8QeUyVY8vFRg2pB8WJIhD3YSPPGP8C3xWgT359h1Y5PopP1Q6PyDvWE/XCsp9DXgITRDQKbp
x6RpnI+sO2ErB6Yn/JZVQTfc9ogASpygTpuZI6kUEcm1aGBU9mHzfCKb4lSTsrBAsCr+SITmViT/
cKvrbn24RNgR8ex52fwaOXl4FQJlh2qTQb0VpYr/1LO5CEr4dT2s26RuBp50ndBXgUH/1W05Fdzk
jV5jxjbnNipVuRYRVpTgGqnS2gpgsSZd8xQbrs9A/GEzO4KH0hbh3bJLMrPH7anO3wv2uafHbPyT
/F9P4W6AISz0XtqEgcA43dg/IbnvSZlGnxJpb8J0bWLyODwMF1wmfT+fZitg+fJhmdd+WUIYSGaB
zyQConcWUblflPvo3muWnTc/618AqN82snlhfHlgG0KVsM2yJybSStZsTM6DJSWepd9WBgQsZfg+
PBn2TcKYJhv5A87SxnskpySl2ZwbSnYJSoymJzx79Rt7quejLg7d/ElHsQ9/IPEcf/oudMJX/3xF
dSS7gVb41qJGXK3BamdzGuam7eaVeyvP1UeirvegsrcUejvyqk4SNKvWmLvV33vIHMjwKR4WcVlc
ObHfWLLk/olHxpRgFW5hs9UE9E8IOKBHKy4nnWrwjU/nzvVCSh5Waia6EJnb1dlN0nivcVN3bkXL
CeVDRiqoH/bqONgGQUjOpNEfuaiDktpVxjBc6fvVDWwQkYrDWNeS+TXWGYyVc9vziJYEC5pQjzkr
vbS9ZauyujVOASqarQD4JKP8T9DshywggKlQchqxk6u9CE7w5fIfas9LDQf8lLysgkAbF/hkm4iF
epz5w+XkPcvA3LTEEPMxKEvliVwTOq/pDpJeE1RsNLU3Gs081LcpvtgRt3jWTzYWw24DDSzS2cqp
B7Z59bJBnW7Z3QzRXAvqjEDI0MOuFJ6l16pUfDJUH33Ux4NYB9BgDlShMOA2POQkMvdk4u8A7Jcm
l7hHccMJ9vUm2VrNfP+L8cuHwbXMksfau41+GsePtA5eA8rKf6sfpVI57Id3mUEgX+5IocfMCsnh
TISQ/R16pOobC8C37nhUeh8K5K6EPD0FJmmy0jj0CeVJ5uXXDAyaQHvxfWTehNUQdeAJLT2vdDPs
DV/M25liGbfR3qfr5TEpOxyd9e4+6NPC7YbYgU4kX/8yzIt4K7hwOVDGP0R3EByb0Ra8YCNQLGKj
wV+/51bQITLT39K3uOzFZzUA3HQow0J++6HdfKwha8/IIjAz+Y2Srlz58G6fPl/9JrbQwpvipW2r
qVvlBF5MQG23ISboY7jYzB1aLUhxg/ZbI2BsadIn2zbVqIAfxisxhhG45O+pnfaMfgjHgq8/s8/K
UgpYJFfKGddFC6O+jdZaa3IqMWFks2bNJHsSm+YNoq3ev+pXRZln0sg6bLF9BPKD+jr9yLvyk4BW
FcoFD/pEXDCJ3TlZT9vXjqd0ROTku41nzRbfjtmE74Ck7zd3al2WMuiG5CX7GBVsGxwJDbttgJrl
J/ZGtPBjP+TK4X4AZvkE6GfS1eJQTz7M7MqXLV4dH9y6Z5ydmMDOsWYx6MYsHU6x652VbNazrsfw
8NQUdnck8ep4Nd+qPf6XwTV6QMiSfhfzYP4plA0kWl/IEITSTvfiSuylF7WC7L3U8s/l+hJk8ND2
kK2TYJF8EXdeRz4lJ9oSMDNhPhCqCdlHnkoYVDLOfoSG6HOvMGZdL43tbS8rz0F6wrGRjEnuYHmm
KMMd9I+dc1N5hIFPyzqkxtNIvP/IGS1t32PClyp94lcx7fgaRBeOWWth7VKji+uNvPjp5wMNYcWj
NqKLpW7V01Dk/0UUig5Xz6WH6bQmEKfoPq5fRZksfCQwsbWLqQcvESUn52a1x+RLLk9ZkIz16bpQ
fT4QdgKC+V5FpUjy4ZSk12lx+R4N2ciohc93Gm/rPh6hd+kyRCB1YQf/SEo5XLiB92vxcVXSrrNt
emMpP4mWNYDHYQPiHC6FuSNi+SNg4OD0nGJNngMN6Fo7VwGVqO4OqtyQ5bH9y0OU1ILx3tYSCX9o
ux0iWQ8Mzp1KxIJuUl/vkQUX/qGoPgxLYi0qc2xWA2jpLddtpXEfocT3ye3GY4ruttrmOD5Ha6O+
TVIgutKfsQVb2N1dKDx4U5KzBkSWm7/mXnRbiF/GMi0pS0eyAN2X1PdnzGJANtkVrWNbYv1DT4tx
viDxUcvgWIsjg9TQO/9DxAPHk7DjWjYv5ldE4IZTp1u5LKVO3Y/efoOIeidfhtudB/nlOvaxb8De
5iIqkmGfziBLWOt1rjokpw6isZY6J3mHkC4VGYrYCIyPYCcmxFe7kTPvHHtTW5usBbZEQDU8Nqtp
gzDQ5fzPu9kERlnXztL42GfLE0i45EFchiFrs9Zn0YfIvP7Rbldy2NABj06bd16Cl0BTM35X2PzO
NPCUHcyju3+Ijb4uIYZ5D8tuE4746z3bzwsUevu+jY4mn4M4EM2msHGXUkojgLG2Rlq/2fe2ofqK
QBlzC1kKan0CHNp0KblIIsIiusyBqCly1YV3IFclNBiMGUL9TBYGy27JtsjLcPwU99AVBMmGdhZr
mGYuIFsaJ0TLC67c05IYq8Fii2+Ji84djksdCvlsWQuSg74KmPy8Z+V+Xqt2sP8N3CW5JkFpK7uA
6E7mLwQTLGSRQicDltf4RQsX6/eNqUSmC2mnljbmmZmMLTCLNwiDUiwtCl2U+H4u8whe9nmmjEIW
c7tleURBqqQEI5rrCTRf2o8H1MZpaPHVVWhVAUx6tkEgtuz7cWKT6uVXrl/Tb2uyIMC2kf0BKAxu
0wyEa30bpM893zS9FboZz66o1+U2e3V/zPToUFMZ/i/RFKqVrRv5cI+nDsGGoHiMA55WaXDctL1j
rxXb2VZSgL23WgHAfTr6ojIf5hawbNzw5ssaSTowZ3n6f1//NRs9nzUbf7BKVgzSDuVEmeLecnyU
MpOTkgdtYl4QHahomybpbmE4kjIo4SMsTDBJnuOk6g+cyLFfiKPypdl9YgUD5KtDyOM8QzsvGTNd
fobL5ym2iLuyMIddJqP79hV8MLJG5yE6oyU0hExMYb6xzhihGjyyvLRQm/sSWmDcsafgEHNDX3to
MsOoGwMjcYID9Un/VkXxFBOfVBCWJms3l9u2SWMPs74vYI0lLBLHKtlCkmV//MLKlNBDAd+92lBf
thp4I5jNJyY1BzdHGYPZJburHmPUsYdQD93bUp2iymb0sI8vYVvYqtBqdNcs4heJHLXg5HZw5BiH
Kn9kMNzjp5GdXSIHh2R9xPLUK6jmQf0DLiLoUNkm5tdAMt38Zx3BnZPObqNy8ON2E3lrpYCAhqzr
AjRl5kvAqFmwxiU6LoICpkrOyxa6LvRlWyaI85zzDn9VWm/lrknm/eGvd2fFwlbAs+NNoxYh4KvM
nZ/N4UkDIcfGtP9E8tN9jKpww5fIADtW6j0A+8UlK2/3Okwb6UNN/hXvqDjLBMYPqVoNtE5s9GJw
MebfuQQ010y15dUY5e6zeLhL/oCb2tjTkaQ+/kE+2TiEZnas12xykgNcm4idpcCqob6znSTntPN3
X9BBx0kJWobbW6bwATIxpoJn49Ah02C5DL5ZRDcGtebjVRuL5TVVgQkQJmh12jbQTAqrmNCrc1ZZ
S8+wCywbUMa90PD8IFG4ZcDddHkOnZBCwwCK6XFR1Vqmduhgo11hdQWmyicT1zLYdpmcj2p8XjQJ
QXZIDyTyNenQu0DU5myPd+t7nPlnAKtfWUOlgF8TnuPd5bKzuMkwkSH5fWOK6LDh7K/ku7Y9UJeJ
mx/aZ8JFdH671Ixz4/3/9tsjAHqg5RnMyN1OrX+v6/fBQHJARGTb6JAVxtoXd484BwHkS8dPuWHG
hQvuemGPlAx8XZo0ob4wJiIDCaWLl7DcfGB/QFPqp7K2radtocOsjyi4bWO1FND3kWUZHsau2kPl
Okv106olu70oGO+F75qBqIi8Hhh1L7ZtYL6V2bvk0y0KDeIQCyuxg4EoVvitGg2s5cD8nhsfG6oM
n2+x/by8eHI4vgIjt+8dRyDGwGkRR/xMqRDlLciBMoRdh0g9THITG8cS+oj1RB+zfaW59eD0wIUi
ELiPrCwRVVINdkmtNPZiziTX8HOM1WyO4DqKKkia/vxxUjbMLVcK7JjskIOFdFuVxLL8FHJA6gag
LOhsElXpPVYWrRTr+Tq2VHB0EqouS4f+fILiUD8nZQeKHs1jaCpYWZ+Tw8Zh8BdwTrNQvbeMtsrQ
M1JBm1GsaRV0tijHrFdVFITrI3OGJrQpTMQoAe6tDKDnJHXQzktnimmXrsozwaTrj9gvpA2NKpu/
0sp7FN3R/gKLdklYR2TKWKbxx0yLw4WBaO1Q5kIuOTPdMGHbbT/+WvCyQg3hy4uSyW1DHfIFYYX8
bJTAVb28eZv827a24FUdbcgFWdjhCoH7C/QWqQZgaG7VHPMazOGr/WKuxDXocZFR6iT4Lt/D+Q29
+K/Px95GiLD6ix/Xub4UiWm8rMSdv8LvstVH4zx7us6wSqc1Ek8DVROONt79rgzbTPshhlIWBN5F
PMAkcrB9JfsbI7HuZMHc+j8TzSD0wO59bBtR9NPpSpPqXF61glE74n24jkIe37YEZk5Z/jW+bj/r
4OGQGZnl1zabvsoY5MYm0X8tQzP0RgtJJDUDf/B8tk/tOAxznslyFgXsnrfB8AlfhacCYqurV34a
Jaj7LnBK9qWqTTYc3BNXODOW1DMBr8QfnBGzYbnqA4MtikiogIKHyCGzeGLQHb/YcQoHZoTiU2eN
6aHLurUN3dF8TkEmYlcTbDi+Y4FJ4FMKnVTvA+MMgoQeS4uQIt+8/B9RNVPlrnf/XWhvde9HToGV
/CZ6J/7WRo4yPzzJmI3nCDJG/rIMRr5zOmHkbOPlwYTHsMW3pu47jnmpIGrsAcgOSjUz63coBIzz
GLCCCRqtBeW7ixNI91H2RLw2PDy3wtQnDluSd3buTdlO1B0Ug9Re/GO5RfUbRvZf1zVIw6ki2tHm
zihYl7cEVitFZ5cvdAHv69FqXyG4ga7C8MUA5szra6U9wf/CDhD+EPvqKGykv5lAnB2QHibh7R5y
4foGMRd3rUkg0ybZ/Mc8nm9MUyFzzvZ28I/aCWWzqmTKk+rGJfoB7pIyhhTXQLKvX/TMPo5Z4t/2
tit2QNePwwGRCKjmxvwOawvFPiLM63dCoIT8VBpoM1+rw/rBNESjzoEwzhMbRAfbF4PNXmV7O6c2
3x5sHgmXxBVvBHXGazJ5gTJf+D2mue759XQKjkLSaJeMDglDoocue3U//h0fbhefHA5tQmst1DqL
N9G2iV+POKJ9oKDOGg+iLxcvD53eYp5Dbxr5TeLx5omPBn2aU5rg62xQCW3UrRyL3RmNRFxYpb4N
bG9euszjBFHkL749AA5uwjLQmG5Sypz0To2MfbkeYTDWfiXuW5jat4JSoDylj1fr6wPQwiWYW1bZ
p+km7Baf+jl/4euF3Gg6g08LzOLyAQ6bfqRSZV/oc69eFVP7rmPCIwVWNGNXl9usVSIOnKPAGUsS
QVTJsQgJh4tHXQO2xc+yw7moQIpSgyvyvHZzW17119w/wGQQJkUg3uNmJ6ZCjhhWDHHKYKhGqxGN
gjM+KgrQBhU4+6wIJksFFB+frwEcJCRihvB6A14Jwq5/PJL/BrakieQEbpYeGBkx2AW5n8YY6w51
swa0UM9778/U4nis2od8K/R/0rf5KeucexmM19r2OM5ha+uZElVeMhTVnMzAA4sVerSBdKaLIMWq
/iNvxdZ6Rds7Fje0pxWQguRkF1bUaPOvO4vturuqrdGAKg67s8UiKbRP3BAviWrE8J3GIDwjiSqs
KBaFYBSqMi1hImg/i+Dpn1odEyIPjACu04DCPrIHEBVBr6h678bFo63XkDIXVC3PB8Z6LtxpBihT
M8McBwn8UAHa7BMZpM+0pSFiYadMi9H9SLutRUP4uXy3KNd/PJ5hFXRl7iviSWz+wLN8n2jIoRBE
2N5gnUaU/dzh+ov896kU/nuZKGVl+f/rczsvBmDzqxEEbpUQp+vsJTYBpgoQhT2fkFyRbI8RQ82a
tMLYgG6OCS1bP4FsZiurjzuHEFII8DxbPz7Q3wAYSvPdk0AjRxgsD40iHIFZNg+mFn3IOg3fmusO
mFM51pEbejoQaalIw33DklTZkc7I6WNSstMtzds3nzQDA0/vJ/tvvLZ8r5Q7LgCA41zRbFTxJWUs
8mGCMsEfJ23v8rpiZENxk+o0kj4pPa42HbumeBpIc3w7RiFmdZcsFS0DPS43PeKiXvcMxs1T7ubj
nFnUYsehMsYzYFAhZjip++v4UMTkw8S5Yd19WnlCeQMKSRdPBuYbdagTgT93gAQhFEXeyMbn6gPb
7t1Jx7rDhPm4ldHxQtPKKyJBAB/jjnIGwXUZiCUJiJCKdS1Ce95Wf5TfG3/trq7Ga3BZ6snmX4sZ
pdsJQJA6hUnYG6V6A9YVyc/cd5MmCF2GXFMqqonh+2Zj4dtXQCXvHgEPi55zuVH6diEwyc1HSYcb
iX13uFR2hrlzyzZUjLOfpIYtD06jzdbLpxeIyvp3L0907DLytAj/lUnU1YITEVtaqmMlOcuOLJeq
04ECs54Yi+d2fPFIMaoygfT7TTC4qKwAyFRip01LsD+AiBiu4jahgAhSCX4qXj0Ymlg5FBnmj/nQ
wBvpg5MSLxIvsqU3LxiODAiUTL6WVECIS8bDHeoVYkLAoSFAcgvLTzmU3XVuz8pF/ibT+45RawGJ
b3HEPJRBcmOG9Hna9SVrkRqj97HTgM6G+eW5MYI/yeIoGnutGWTsco5RsBrvqqu6njr7ERmi3IcI
9/BDgHpa6CTzUptK5qrsRUHtMqaB0z/x8asKxwcf3X7NskhIXeKGND0PxVM478LDJ7xckFrez28O
EGe9lYJM7zBqR3oldDzpv4izoRbSwpTQxvSz1Jcx6DISmiIXuQdTp/qGvQ8iAQXA7AtSXpVxmnvf
+U0Lo/GRb5uthqyppQZKLzwOoIL02HYE6ryyvrjaXtdTwNJTJi0KzRPmFSG1y96QQgaEHCJPLFVY
Iz4LaXjDY28WUIblaJ3nEsxLHxUV7PXX1KzkQ3xV57s4JR9l+E24LC46yECICsNhBTtE/FKDWqu3
oCDAWHag/oWR87+wAlnXhrGHDB+3REyvEjEYnR+4lfQ4CtzjYMEj1VeiW5eA6qjjxpsp9dHS0cec
u4MPil38Min63G/MCxXiqigKiuJxaxej800nRcFCg0Ppm/yLXXKeH3eZ1Ua/bSr0dmJYaJUIIEf+
r9ZQLTKrL8vNyKdcq9Z1y4h+JWrBWgj4yrLizDpJAlQsmd6DKg+L/MzxssZS9bJsJtVMrz2c3cSX
OS+GLvX4QPEsbDIil6SKvTFppia8AKuerpQIpdbIXulajP8JaJFdIcSyzi2ahlSecpprk+D3G9pa
Lcl5kqVNflBk4GuZ5SKYIJenqwXGclLyUQhUgeR1kDUG+n66qZ7d+HR0Cg2YfC060TscbxkuXClS
xnNwE7/xp9fGgVlJ0XMmpB2sWy0Mxl+Z6kSgiHqP7L7Afc0rlL7lebQSQNf0kJCyLSDxB3nphI17
evInIe8557elEb3cXcpTm4DZtKc92jwmYob5XxDy5IkaB5RMz6GZXKxQJ6RhorCF10UC2Wdyjl/e
wOKmnRNBaY9J5R+kU35AUHz0F+PLLzDrcj8Eju1g4/HgEs/1yZEGlfYtCfMemCgYMBtTtqnqihQY
Up4/pa0AUJ+PFE3Tlb12sjDASRGQLQkW4IK0MbC84sWb569nNRCn5kzmvcLlS2MR9BDoBXZu5x7f
kaghfabyfSFGou0LgkuvADT9vrEEeOk3HfmyhI1C9UWUjontssEBbeklBWf+1s+1iW28asq/+vgZ
nLSkWG7lE1roFgffsUe2EwyDhmm+A8IYvJAdn8taYOSc664dq4a6Du0zMlQkugHE11i2Be9J3+fE
/BY6xaoDVOEG9GMLUD5F2TYAVXt52d7Y/yB2c9IFKlTxlaB+jOqb9IacifXymFRCo0SfIZ10o0ZS
GqMjRscsE6PFWh8Cxr6Z4y5GwFVj0jv4uQTG4XtArIu+hOtv93kQu1aHadN5kmKsze7r7PaGdZgF
F0PqX4pYPYewyuty/Y3108Qdzkz7HQ9AKJDR6q+pCzlzYHieNUlRd748PQh6s8fmn1wf/ECOV6/O
dvJc8GH8mCwa0S6q2YT5nVteQraOBR6a+Td/wscdXLU0dmb4RuW/Fe5y/zxmn6HUBDsWQGXHRkL0
pADw2GtNcz7ahUwvE61gZwlTO4pgaPJklNjgavxxo4FBW484jYTn5zVH3aRWh4vaRHPFHodV5XnS
ZypIfPLRffgZ01kswJfNbDCVTuynyk1cvcEHoqHduNDrQ6m8gVl0EnHNcqTDjWs7ZuoEA1LYFjze
9xiPUs6Fq/YikiD7tGtWN6bMQb3/NzcQxWy/p3cra7yC7xllMOEf5aT9wMOppvA9R+lQEmAFHUSV
IB7hnmnO3HJokNfHfqe6nwe3FZcXRppGE8l8hZNIHWRUXN5yHOljSjZuSwY46ltVPDPfo9xEP4w5
bKRk6SiEGMp18CY7U8J/y0KjU7LR1bCBKlbfIwXqueL5Q9NF+SkaVVV3eQqmuHj9lupEa5KFG0N1
VCttcv11ZqTdJ32mIXKEO9l3S1d16CUJW40kotv9s0YgzJiPCPH5qNy34GXbuTr1N+Xz2cGUSQK1
4xVautgmtjmQqMpCrl2ckIXnSvil0jXl3HBMVeXvwQJ/OTUAD0hnSxVBxLuxGI09Y/8Gq/rGSM9o
necVFDCMnEaRa93vk6D7wqYU4atvxYTcxry28zD0Q+uXTFFxkDkEeR8Vx2KALnbFeSFpnalMbisW
oihB5r9yQLuzdhdjpABXB9KUUbL/0lm1vCSHvE44nP9nhEiGNnKZ5fFWIZddX1U33MbhAiLohxe3
sf0bv4iPSQOWDerU6iBPhU3l8jexOeirvHBhLlNHshaDOLe4dF10ip3XBX/fdZyppE9ibmHYuUTP
YbWzqIG4kw9YrACPkdQ7YpI3VjDYVhVPuvyQlHyXBcdiSpJw3locY2yIx9x5utXks+0AsJONRaZo
dF7VEcPDctkG1DDURmug00peXfA2QHWW+NzHfiB3MAiwageEs9QF13L8Jo296QUhPJzjyXuuPr0W
G7/AEluJalaChyYDeMfOV2CHETdbGD9CECG/KmHfwk43r65EpKI+iS49Trs4KkoznrUwE/u6fn86
ph8MlpMJjxG2Ijp2HVPZtKD1X7/C9KXK1+ztv8ppelmTNo5jXAsYjEZfvTkdsqFX5rr3+j4X2dP2
2gAR4e+neumcH3zPKzdUG+OThTVI60eF/pHCZhJH5oXa/8DifWg7CmfGJiwVpG7SqItShJpaB1hS
qnaazVsanTe8rnBzvKo9oCBmj96EzWxLBEnf0zm+TzvzcSPMxzxhxIuCX1JvBsa5qaLEjj3LEeGS
DPpS4Dt/jO2exl8mVSFFvAQjeqrJWkQ+IZy98teM4ntAa5i48Vb7w98Zs9PrAu5ckEAJ3c7JSjTp
Fj6M87a6nzF9rPe1mxsh48eDt1p6trUH3NI9GB5fXXYtYRxGrtriehzdKdSQ3yiHo/cAVAKaoOqQ
8ilzg8iuFrY0DC0TXyIDRISB2TXOCzDkE7ZQ/qcZrUi095tn6TvnJSjhfiRbm1+R6CUKtbggcBfZ
VinhdUIA6KOTagVymOLFi5jFJ2wtYM2PvuSYHxzoSNV9h/NEKBPut1TxmpnlrQ6dLIqm9tMbFlGt
OUcA7uqYDBQR2q6DuDkLEuY59pEXs5z/OatDfVfg8+FVgR5+8R2/suUpFeuL1zcP4Acyq8FHFwI2
bmQKHGNcqYc0Y6U4BD4/qarJChjIFNc3f88ZVZzTR2tskPihANB4hfyas4a52ub6jS5rmBD0vh7l
XgMbnIFmkqhbv0gLJwdql38qahtIwJ5pz/BeSeC5dL0U/AdZDtHX9qF9i8L+K9rNrvdSfMzEtFfX
OGuGMAWlF0IQuy17dvQX63WUzGCBvu7G227iMouHtynJHiA09s7Eor0lYA4lUd1Rgk4/LC5vm0ft
NzgpPyAT7y59Bh0A+ui1+J8yXWDi4Z7cXXZZdS1WTyEhk4nLksmn56NFE4ZNf2PHJS3yHgRoYv0X
5pIwxZzC7aUSgCMksH7zrkFcumlXvD/lhHr4MY0vnFAW7Or4/yAbt5zKAh5ZNE7zk0etrIoav7zn
daMm8t1/yXsEAJ9kLgmOXDbJa/TJNVxiPXtKGgymkcJTIC8ysntlFwScxlWW/RQg1YjLgDqgQ4Zx
IQxmMMa2wUo4IEFmos/ZiTmlSi02T3HzFLoaPYZeU5d4BE4ajfo5ybsJTUKdcw72SmdwyI7jMVoS
XsspPmDWkHJgJEyoYrnE+SNW2IZGtwCrEVVT5X63HmXQwwDLA8F+/LQlRRXZtLSRRb7kMcW275BO
o//QDb3gbfbjZlbndKwCzP4K0Y20LIP6QdeGLqIAf/AKHr78rP5diADNRINhukEy5OkRwWScjfUw
3qM6uUShKm/i+liPEJcW8ezVEkBffN/WpN00MD7iZiuBsBTVdYo60iuQCexU25NN5CuKVyaflo1K
Qq7z1lPZLqZSmXmqOaA/M3ytgH7mgXBVx/GkyCNBb25lbv90NIHrq+Gd8AtCE3FlHCnBRx/+CVwz
aal1vDQCMZnw4knVhMyfiKd2EaKIjksDpRRAKrNzocklY54qQUBHCZbIMtBS9HOsu5BiuvQWdiMn
NxEpDzZYsym7bc5W+F39Sr8DFbxN0//GumeUMuDyR8mNbWAlrhUFsiO5KtNyMXSmRozJ9Qu5UGup
N9EdwsZ3+ebVtJVq0nhxFco71lXJW3KHgvAREtYOcU32OkpLNEjjLL85jwWKQ5akUwxfzdkntAnd
U4iuMVD7uEtHxyqwK32Q684/83j3rOi0FSf1qbwJvy93fH/UYN0dl/7otyIzzHG+zvO9HDhS3PfL
9DwnY5uxoDXhwNgJY71Cq/VcdEkuqFLG3Vaoi7kqzFBpzgsBgWC6oGe9Apgd8N5GIStcAPgoo9+l
XD/CPteQcn1SOlCHFgRPY96458kYYPYT02D7oQN4eXIgAU/BzJLgi8mCUF+DhnGdgNtoyfzydeIg
+lXc+12dZU18SoyhuTQqPg4/O2sAiH9yNaz5JkquDmCR4idNalO14fp/I1PFL67Vl+Xa3dMuwDg6
J2biUSfhFtUaS7Bwfi+LBU7tjPv3VjFNyuejHJ5xLamRocTXPThwwDctyQEORe/XnbZCEQtveTVT
V01YIoG/SPbXalPzBCjBs3Ty22T0dtj7cTMuOaW2LtyZgdT+cmZMeGeiY7s1LpmYvjUytIk4Rvhh
OuHLHJGRQISGOoCXrEMHyc4zGO4l99pOlz68zlGir3tDMI/crGCKgQcV3gIeyrMHkqybAnTsM7Qq
NPyLei99gAtSy3sYVF4j3xoEeQo46Fld4BmTKmHqyDESqcFt7gIsmStBq19/ZPw97Py7QyoWEo7y
eM3YUqH3Pb2YsorNDqoCkPaggTiWLHnNETJuKXj2+tAjrp3G6O61J9/mlvOLL4vyuZb7A9AGAxbZ
KTT9JlK/kR8PcCCvc4M9lANOjaao0AEpl7YnLKxEW6vmdGM0Xq86Jmmuel5SiEoqmXN7nJGTrzWx
ptOMYBDOsOhbJzYEYLCK01GNr1/4JGHFFJyWyer7IpIQsJmtVtK9frXAJCQZ/qjD9SUlzJog7A+8
Yjuv1SYLaTTJyuBfXRxamOBpTyhgCocByluSZ0QSv7eNeTqAJiYvCPYH2ZCu4EQ0tk/YaRJRIQyS
3zsd7LjMzJzKXzno1BswHRzepNvWA/NElwTY1vjZhv3j2k/oUdmWSM13MTBybAoeQHZb0g1Hk/tH
b8BBWq5RRqw67RvXmerMxJ0q9gX3knIaEiDTnkMsIFsoEtPLL0f+Mh8uaPsG296a4n6bjB8Qe4jl
Y82s8XkOgZckP6Lsl5gkFyEhbaI5JUKpvNX6nbVfFmpmsc3aR3BdckkmHDUS4CC6VodYC9j0x+W6
O7SyyGVLjLPJz8IxzVoqApH+N4HLTPsqeSut0MjhNxOXRxamMsQfNaL4JLbz9Dfo+DbrxLcP97Gy
lyE9SQVBQfH4uqvwTH4LduvAqQZSsOgFI6U6FaKsTomQ8mtEAhoDyaM2rCw+BeZXlHb3c+AZzmui
eqmk89qVztaEeLpvmWtWwvW4/eBLDWNRcBbhvQWUggY4PCtUtBixrJK8e9p/7DO5uBsca8fxXrds
rhtCa3dIwD4AH/9pMxbTiHKCRnMbGmu4b0HYTv7SLjGbJOIadxyrejU1x0MhsejRPVufCK6QdU57
b+q7i7PUFVy3mNgHkT2wqeKTT+FssZM57dIeWHJei91ghykIiFL5VrBV/d1kCo8dPWgtxaYdlRsy
GM05p2FcT0SosNRtVIUmM6JEnV99bic1HsUvX2vRL8PT83mBbrRv1zm1QCvv01G2T87oApKlA0Cv
ZUab9i9FllPEyV04Ok45EyBhauxju2wQg4VDTn/80Z0UeWHFkPk6SoIYUwEJH5DS8s9HC52SSrDa
lmvxLaoh3cEf4dxnE95FCpkcPo3q/EgoTCzBSUOaNb+KR5DsSZdg/hTCvcmfbdhnpPBcq9WA0jma
2UtloqxXFJvnUsZuIGxl/xMI7kXGSmrOFnNf0ZpQTzDgSUbuxMQ6A6ifkwNQBUpG4hwDbEQtCYE0
q59XUaLstB5tylxC+WK0UWyyR8UlOX/yCD+oayIF06+W37r5JVrSWHT7viYHNdotRzXUSCMLYblJ
cwO73xHykOTcLoqitiOk1mTOihED16Xy3Oi0c6wi02T517iQdGjg8pdevNYjFKWjNDt65CmYSHh1
lpDZQ4XohPjDM+KZHiLGYKEBuE8BfXK/E+cDf0qb66lssrsbztRt/wGE2luaYNmtUF4iwO/t9itW
McMpC35PHYLejoe2DnoNivcqA5zk54Wg2x04clil+LcxLLXOaKuLq1KAd9qooyUSRmH2x+QE88iP
trM1Tg9uUsVAnQAR96O1owa66lkXL4fLAX6KAwgvsdj9V8yhZOHmcsYWqTWb5LPwnwAessRQjtoO
4JzkPuIyDdYJbsOjw9mdMkypmRQUBr7hxjey24axzX9qz36sMUjKa1t2x6tHmGJvTqBgipR9XSE8
lWGd7tw/u+Izl+l8KxKt8ECouFowWjZE35I9oMu78lTblznxo2lfyaX88lGjCdOMhLLzFJtmcylq
+C6kHkRUdxUGDmIZvx0kpiAQdU2okHoBgMFpuUP3BT1aFdFxtSFRaXKGICi8Hf48+YJ7a6DIH4jR
kwdRRtBW2WHF/1OIz8zLk4sQ4S+kb9RYARgKjIBzTcO2YF4G/KxVfa4fIxYIPpy/zp9B+A0M78Ff
wH8HYKb/OsvlqBy9bC6xjPOB7+RpqQCDd9/AXYZ2mo+o5C/UzrRJTzLu009400pcNOhvpKlrb7nZ
EyRIMP7JK3/lZJsY+y8ArbpBCW7mJenQjlvGobUOOq7ulNm12ZbWcL5UBrdejqmpVXV7KatBcXy/
dCYaBtX2f19uibsisIoThv3wfdyUu5NDcmnxpXRWW/qRDurVfb8JmDheeNGg8YMil7k64V5mb0Lt
uhHiM7Hw4H3EQVXUHj9WqSvH0tPllyBxM0c6XUDPyDTBQlQm+ykFDCjMiqO2NkMUdfFKmpkTqSb8
LWsutNDOGD//l8Iq0NASHB4KwfwvW9nMO7bnBT+4ph9EtNp3i+eciXXdf6CkmcbQsDlFvrO3beSA
5ADisWAwxjgwNUu8LgsWochXEYheOI5g8mjMoPku+NhK8k2rrvdIYGx9mCiURioAAKLbh6yJLsnh
PMTKca0Pb3I8rHUkphOQT9dTv5L35QEEWTSE+mVpJ+xUouT/LOCvwz6VZFl61hoMb3tsszRwftAX
tvNlwr0QygADrn2rUJUxz4uwKGesP2wux70MX5rL+zcXco3Il3L+9m0DhA8fqe+EMVPE4TmPOYrU
d2iPoU+SjFA3fryHgEdHnsmaQbD3EvmW6AlrmBWYjJbAB0vIgSeSQBpFCAHgytWRU3bB1SOxMgau
Tp793yc+oNwlFBO7KZeFPgM6ryopq5CD0Yq6Vm6J5omceLbpkoH+RFPcxYbtg16illLb2esvtfd2
6LNXWUf1B2FuW/nvnBw2c9EWCczc2Ps41TvZATLvhV5jTuncX83AVV/t4Ln+lKWsF2Q+NRvE96k/
v0NS/dhkXktwhzfkwOJxvld9Nzh9V/CiiPx2E+5Eh8E1RDupB3Rku/9FLWIWU/5Tvl3iEF9myp7e
nEh7SdFoJhHW2anJ+6y7y+m7vQY6LUFHD2IRZyIBxU8Ro4k+kqYUprmR7LrTHRA4UOgoqf9E7h9f
GSEEVDl/vR7Is+1/Gd1e2i+iKS/UNDBsYgl8sVnmj516UVDJFVlYc+2eBMz3kM5EKSCfYUp9yToo
FDikA7ys0OHB+xOJ+jY8gOAaZVdlSz+1way7fZBv18jSgkEwchQ5mTB8SV12g658EHKz0EsoMh7H
ui/kb1Nnne4BCbnqrP688siMuIWHO2eL7jqyyiyU0e+8TqA8Rppb8wnO7VJWJT8Q3rUdXM/yZLdH
kZRF7k3Fvnfp6ISFh9AX61HjvvP3hEAuufZu1zDRpPp6Wx7EU6K4B01cShRa8MbAG+KpOwSSB5qE
7yg5ttmtu0B2+xoIuPcUqkUqE6eBZtU0TXJ9bCduo+acAW/oQYRrRWiVUZq1Avpkn7Cxf1N2qRYH
GCQyf/6R8dbT2WrR9pyDGx6mJoI8fum/J23AF7ZVT4OMrDD7bRURo83nFXIYtL/eEeK98jaKMahc
FRFR7Vc3m/iI0FaO7RytL95Sq2TlSAMKDcNpRmwbifisVWLZBzhA7rZwWml8Z0JH078/IPglSdcR
0M7XfAwtQB8ox8c5zNC948Dk3T/AIDlmPcqnrfTMMLUhUILGC6hB1e1tOAJ8pIGwToaIdkLp+BMh
ZBKbepV4jrbv7PD0eYL5f7xszng+tWFcebtYLQDTC4xtFX20CRDIh1FDVMwFEeH1Gu2wkXy4qIwl
ul1Ws2+dfW2qIg/ujJuGgpEtNhmaVdiYkb12wxyqzOWFTrSvNPAc1OqM9Q7yIutVTv8FcWaAEu5Z
r6DGa18Q4vv2kL/7zaQzG3hk958aMNmmne1pBZ/SlvKrfacaSyAJ4qhqnSkJIkBP1ZVO6WPTBRCR
zyiyHJXZsV5eYmWaqz0FL9HugtavJiAbmwFSLy+MWaT5Mig88Xfj1TTwhsiweGrV1fC2fqq14q//
YX65g8Bwq5FIagV/kLNM/2vlT0h96oxZDNiZasYrBZboUFchLXL5F+aF5bYkOXNTvLLK5dTlp/bR
erQQqFBu60BP1ycW/m9+5W39xmA1IJgLBS/W8W2XqUrDtbeJJN/oZ0A4XG78ZXzrk7BrWiBq8HVI
EDUSHbH1lpgINGrWd5FLu5FGbO+M1TgYNUtuJpBQ4lg6OxNYki5dsXAjSYDkFI1d9E8OLRu+MRgV
LW+YCvpNfWDWRkkyLOAEclWTcQe2UsNx4iezf7Oov7lRfKoSF3pqMLja/ymRiXDPeNvQ3mhyKf77
L7UpO2+3bLe3vBBBT9oorF1BKWc90rfbSNtDWUPlIwdSyczijWH5WtxG6GEpBFqnPmlw9ZlZj+pa
VjEafiD8aAlIZq0ojFsxQxJidN9DOrRz//BU+skrOygje9Ddzvb1jThyL1SFoM9bStXVon9uOXvk
FcB95YWMxBJ4xlhEM0IL5eSj1KNxgZ/FKKXpOvLm5QxcaOcj3/sVFjoq2re3/1mnWWsZaxFiRHaA
nlshlMGlYYM42AlgoIFWhlx/nKGIgFW4lxQuySLMIZtTIdSxf1rpUSCU++GfiGWuLYFW4y8esjun
KrGnoWIVtLEDHXwSaWDx4kHHp2ZpGAqrDDJOo6T7BMv9ViqZzFvMHqmwhU6e+JILM+EFVbuj5Y/b
MlnGRk2F0vdiZieUe3RHb+JAlhR8xVz5S9g+lZdttfGgL7mG23qae8Qczet/0tQRuC6+MAKaXOkw
t9Fr/VPbN0Jvf5nsPSS4AxJCHliVlvveBbL0Kj62YUISTYQ/70bZmroZ8x7nrYX7ilNePGathxYn
lu8k3t7xWD3d1w+QyBuTkqBIjNN75W+u5stlyr3uTtiurSmAma0PtCW+nijs4Dk+ovyp5m93JHyM
t3ZW016pwNEWeS+rvlRxHSI71Ybvr8EjEIqtsrDJRnq4sIeXhYVZ7GPHl9ORGyOQUy8mL6Ho7DMx
FkbJTcYZPoEmJWtIgiZp+Cc+dpi00qSLR9/rhtkNTm6iW5GidRyXWqS4jD59amEFSficlt4FmXT1
NkO5/b5tDnKffG/fAnfv2BaUVhu2t4PJujlhRoyg4X5nTjEtS6+87g1DYkwe0YqigP+bWIdZsdt0
IMlAt4/LofF0Lk3LQ7fqaAPhbsrkKOoLLKryUXs2QUtugukIbhFhYg5bSf8i2EecV/e1ZrJ9KuYz
qnzQ9LBHbyvnQtYmnsC9GQos3WFs+6j+HFVCMshM4NKuyVMI47ZvC8zYokm0BZhwGgHJ/Xo9D4Ed
29oKu63Vsn8JR0IYmT+G/8PiB1eecrasfJNVunH9Zboke8aBi5jg8hWGJv8bbQ0mUgt0Lel9shYX
uZf2yjsoCa7D1PilHYk9mvIdS/9uZfxRUL39RZTr756esU2RGkPwhtV5YfOvzOWIuT6P97vS1bE4
GBRmO7XL2j1wd089NUrlPL0VFLHLZWWAu0XCanXaRgqZJt9hLZexShDNSiDMdhpi6dd8cTPWdDbA
Nf32OWEIozSEMfktj1wyIn47ObsMPB4vO7YoMzND3ZWi/GBrsjoIJV/s4hZUf+FVigPEpZ9enGJr
hxntqmPzUkPJLTlyaKver0KJ58Hvsf9BBhWV/UtwQlZGuIHklYOfY/BT7nHaT9uQfGWBU1IXJyaB
HFbhE9Sg/pppDnFRqvlQUuapu9bu8qLRLIAgbvk78DWtPeorsDR1IAnTMUyzYCNE1ywmUf1G5Oam
rgP071wSLfdDNGeYJPd/lMvVmN6Cq1MeZ7rXGwl1SXZJDana/D30WhMxpo6nNqZBY/ZDa7etEdMf
98M3hnj6Y/KjFwej36ruruXDs/9MsNnLT2Lwl5HNGz/jX5ZgqbdImL+Wb1Ae7xEfO1JZZJXneInf
rHTRwvzlAsupIQo0U2bVROWOaEP+DqOM8f9rWb7rhUVfwReaTiN4FFwAyNEWFSvZ0UfspvjLR2xb
6BFjN7JJw+jfXgMxdmk/QQ1WXCl2DvhUE8TSqz1CbD08iOzCpRU6EgNIQkGaie0c788hpTwpeZgZ
gvIvoxt4VqU+TLjaAtmC4MjTn2Um1qv6aM1LFdDf8HFrde7wJSOngwQDWWZjAZAd8COCL1ixGZ8N
qqtd2K5sNh7rBYa+/aVNhU514I1ba+7v3sDWcUBw+99y2KIpCFDEJv9gU2fZRQfqYL40gWR27YkT
XuRhRa2y4b80iLBa22wViwCAXFtgIO/y0d5apju9Sp19AYt8Z0XZqjwhtjMdkF2vaIcurPHE+2bN
hVKkkdVvb6Oy4W6kyT0SYMCokutuEmyAdvBevarPNQ2TTBM6XC3gB8nXHDdZ4HrVtDyGT25dlVCY
2YSOXimeiHVUrV6snjgkY7Qdnlw9yzeEtIjJ3YDlgkwQ+ml1nmaWcEBJDoMfu4CGfJbg+J0xsQ+p
rAfEmbj1XYR/uorK+EZNMifp2Ue/Iq5/IgA7hNdspIpX+WIEKooLUyYt+82Mk06AFe3XNYOrmMHp
R9MFlHBVcCO3kmNv+teYntouaFUziD4fciL5BT/k1tLWQYIY5NNnzjAQX4e1sGGtY4bNpgtnv3RQ
HqER/oZ7WCEOQof8NWvPwdTUbBFGt8tJyba5v+09r5cEJWiXteX0XR12VP76s5gziVA4nYPZTslz
LCVd4Q6XQkHD+d6SFk/FNnyiJZHamYrWb8iVuYVT9GXxAVQV4R7a2aqi+YkfVbzSlrtJOxdqlAGg
2gbxPizvWHCxL4gWt7pG9uyvUbh6ER/8hX1Y1N015fG/nXV4uSPi9fbXHsV7lA0gkEQALgRWNufJ
aU3oDCfk/W75ZCArXEYX9Eq2O49zsKsq2bGChdjo+LFnpFVdt9H7pzFszK8nfgW81SviOj9XFwiY
oMl36gpE13FD1mEkyE4/m5VmS+tbBul9+hiPZ/eoYcb+ls7y8XOQFqHAiPfIrPs95x0VQh9sjdC3
pb2a/isyj8soptn7/NbbpSh3lQUY7wzsonPlQVLImgnyEd02DtkgTBFgx2Tvx8hDCDQcR/eHkzrt
EBZC9QGVI7QZ4TGECI7Btg415WrIibJK/3YLbwoUZQmORd+u071DsAvC1AVz+rEPxvUMFyeEl7SP
BeRmtXPS0Bp9rW1RtZZJFK+cDkS2bAePxZe1DGg4w4LeLAS5rw2kF+j2IqvqAwBSkOGqDkRINYaM
DAKMA6v+qf6n+onZCjkS4ujVSK2XPIaeW910xcM2gFtoqQswhie0+OatTVgOeEyHzPeO40ofqSX9
QyZ23l+s6FfkCnYMxgM+5RWIsBr5G4G2Mgs1yS2Mdet6fKQUUpO6QyO4BTD21ZfG1KgPVyQPFpn5
EfPrl+IftX+/DDXwEoL1gbeCco8bfChtx6UMWKMnACNzFFeiPlRovf+tZM8WUdbNuUUkpQ/clkCx
7XJCrJTRQ7xh7sgxwOGPQbz6Xj32vGsc+954zit4FZVQNAylEK+PFZHlYJWgBaL+NPxuJnciLXBc
3cUJvQfVhUoOJ0xRRW1VCtaqehTf+8re1tN6F2Eip20W5I26E3GfL3MqtetNdS2PEuc633ZBlmf/
7d0MS+tZOjywHT3qXi6LFUycYWe2pS0xVb4fUqKPVp5E6on3YkmGY/qsCIurtcw/MoUV9VOblBax
V3+6uaTtF5KTkes6Y0WTN4W2VQ330Z3gB6L5DqUXJEjs2NEUE1rbubaIVtxkPtYYW1l48d7s2/ky
vN6jBbPLSDg1ZgBHtwAhWhf2dQSrQjHv2Ff8cF4N+OCXxbGTb2iLVtBW19q0ONwRkb1BuCDI/7Lg
7nwnInCYVSJfoaZKU9dWgee1GyE0OP1kReMegufe6n57lDz6EVH23/iUmdrdcgm9a8GyhINq/qHo
d+iuHuOeKt+vRlcd2sxaldEjp+zpJQuWZMwlCpRWmI3NfwRZ2sjUwycWlWXfHRMd4ltdNiHw584h
DOfPf2V7nUlj/VAYSQfylnHIwR2epRjtsGRGMCMpyRtAy1JZfGEv0VV0Z/4MlG+Oi/Zw/ns2gnrq
eZSxKMNizdqHNIrUfC+WnlO9XkLtVvPgI5SxAhUPiWXLPUxq0nFvq9dNT78HujbKW/d9FUxfEetb
MO2IOanYuLND7FWD4Gzr5+bMb5+U7udPtyXp7jfVVRVHpjWZ9VJ3jNLaFGjuq+TVw/mTa2KkiEYA
XNtiT0VpjeFkhElAy8tGA3CpDTIZrs/dFteerIsSNGitY5c0gSgBTRQmNOs3NWo9gFar8VbcgvLh
pdkGaDYIXlWB79daKwYIjpqPE1A1Y30DITJ9ddZ2LGJCybF6aVqz4ths6hVtySiFG92esf0TRdUd
yV4q/rdtLeQhWT51mrBtYlPDHMxVDLGt6XM2LYSTnAnr7N/DaXFoshGOdt0DVlCWh+Bnp4/jZSu9
6jRlbk1XLv1wAsFjCoy2mpRTzSpww31cjDlkJYhWjrmGyJ8sYAbs+CCWvpvVfnqVlbTXINU618LK
o0d2LtgqYoMD17dUddHv+fZomj3ShHszloKOYGN6DPkW1f3g/6PtiVsuU1OvlWrnsFlTDJREmzUJ
09G4P8vruTfLSA3YUkb1BqNWeY0x5XP9tbdriiiR4sB5YcZu1BSObMkhNPKQKc+95lLdvAVbK3DD
XChtOAODRouceNbiiWqj8EnEf+N7AEjgUEtndnWYTpa9jxFZRA9vnU6qDRv5B946o6N43glLlsdW
qSgbrUa2bQfCupjqi/aH47dxIBEdZbOw6U5PDblQLAWXzqaeAP3YKCxiRvX2oZ6lzNuxcvs5C5Cb
BHK3tX4gqmxooesaNpMuqsSqOhqgU5DdppRZycm2IJLLNK23S5UHEzMZsg0YSmv6aXWGoU1fOzON
DWbTXxV+IhSktw8oKyFbXA/SEXqvtOK73PvDIftSfeG1K+Fof/6iyJM7YYEDSos1sTRAcz5Fe1rY
NzIKfgv8OsWK1pXMAJ2QizwE3N4Q7nPzf1B/wLPFLaTBQMYZu3Dr2KxMI7J7EVNGnR0gQw3K002K
imYgyyHJlu8qvwRs8I6ToTZau7YuAVkUc6R558QmFsp/9EPkNmEAMDvhmZIGWqbwD6ohiSQ+8eaK
mOzuL+iU3ksDYfBifg8iuWgxTrNI+xTtOxfwX9YtH+HFf9wT4jyjpRAmpn5hoY+hZXgn/T7xXGx0
Q3UiRViGrRmisSV2XOpDm5dQ9W15Ux4wSGXnqqOFHciWVh+kxjfBZW9PIVueqYnFr5FD31KeTNJV
Gm76zubSVDR2RKcyFQnMqO+wX/aSHM3c3ZNVCqEa9PBry2M8tNL46Dza/CtMntg5sUsKdKcVEDOM
2c9mWh3FRLDKbp+y+Klnst6ZLJwv82iF78hRqUFjmXpWOHmBfE/ttAK3euZtw8ccc1nprMVibiQA
Pd2KGWi1Edw4PFcxuLWH+UPv2O/GeTOV+Hj7i91q8aFhIvVxmk6i6JBej0IFGvGz81NXxtZva6Jo
6iQ48m8e2cmHcDfO2KOU89Ckp+5gm4+nXXvGw6CkUXVK+uFW+8CD95bhnWuUE1kkiwoCPlwFmcGc
I4b0xzlEL6znM9EKDmUvW9BxuDDU8fnDvQdbecEtiMOIH8aCEyfEsp2ul1L0TZoOxoepKyyRTtth
Rl+Ivz4vl28FQMPUoUymdC3/J1/4JepzqeUfZZ8o9W6REwajWIyrZ1xLmz6Q8qCpxUgSCbH9bl6r
dZfU/QNKXgbZOFtw60Fpn58mjnqjEmoBrTZJ9hrQmJUKNfhf/j7hSw/sNTGMy51+czKB/iD4c+Tg
vAPbYGucNjIjC8mVsMaRvzIpWcleJKRWF4hBxhWCtRReG7HYdJkboOnHMSXGdKrfKhk3e10FN52Y
by4tK9rte5xHfS/LhtRiyTJk1UgOGksYZwqYlkjatiUYUQAtOE/6LYX0QyL4q4QEkUGiVc0KpEB9
vxVLAydkfYWmCFW4GCAJ9Wnw/dZWz+3HXv5if8CAzEDH5fokzNNa3+JDcAWA+7OQeT3swmV5RFtW
7WscjJ01cNMLeYoEqmTnzOjx/Og6MVWh1P5DkcN7JgCdhu0owq0nstvbA9vQ/YDUBB/yf/9Ap5ZR
6f50zFndRgKCjL2bBHzt7NV+zBCKWB+HoqgvvB9G5o6eTuEcV/iu9zaDYT8C3rguu+6PMCI+g+BG
NJ/AyUXBPpmQODK5iFHSRlvDtpibIFmNUz7wkupt7vpD1evmbwA3OgMYTg1+PU/X9Lu34nHcs7zw
Uq+OcA8Z4T1CAwsnJIQ3r+be65t00ppb5BRZbkpTVhP/7hX1KQcYAFGshmTCmTMC3Xph01N9HF7w
f5FyV/I96OJ51+m78pKY2M6UfpO859zU6RxmfttaNJ/pum4Zfz0VczE1L3b5lbr9+QjRbHt7LJpw
S6D3LBRTmn3l+CZBPEwCEaTLmWcSbdtO4jy3KsEusuhvFeXvz/2mjVyEcYWxggJE8/kYVqQdYXKx
dvDXkuRzA3NrdMkxayjAhgjj3NBI2QjOrjG2TuCnn5a0QJGAY3nMGkLkA7agu8sfd/1W5q+ndYid
1vCcprbVtQhi8evVWbB8myH9elCSOfxyhzqQ50IiasAM3vSN0M61NajVbqA1TvMNH+rkEnCF9Gv9
jZmQwOh4AxCrhsm9ZOyt0Oa92UK63rvLoi+vj54DzQpUMS8h120Z5+ljPHj0t0ZFFUcZhID/ydgH
9EV3MB/wPvod4zohLvV8+r6bMy7RO74SMM/I9aBDu82sVjAWO/5FWxjIeZfrHHAsyTHpAqeywZkq
Ech6HEaghL2nLhPd06Il58aONISsYaDEz3j1SQNnc7nAuNCnTLHED+h1EqKzqcNYa1k4tKw+N0ka
3xUnlEkB5rGUr0Gee4Y+0dRlIip3MpaDF3OlYESaXqGjtNwQP0ASXeOrKUJXFjnMHcI4TdtWET7y
n8mZ9laG7L3B0+K2v8gtcG2WSQmxaX9B6t0xf/ybpA0unReHoluchjvnAMBPijUgyeXjb2X4fzDi
SDBhDMwHYsFXvx/PR1Y7PbD7wTUQIqXMWPXD0eapaNIe3ED8WRjxywzSPlBjYInico1kaEAfjTOA
DTb6bsHhA8iG1IzZp027QsmbihsgphcSJU1jFnrSjVW/zGlDEBsJBD9yD9pStEc64pTS3Hjs3qu7
V1hPEz35K4vnYl5qrfQWlyPTEVyyvyDOFnxAGw9Y282XxMHGe6KC0WZc6Zcn9dK33vOqLJq98IXT
UmZB/k9o8ZhKVvNNxWcKwkvC9mXqctjx96HngztoYk2n4TM5ewJ44KPdO8gvqAWEMJMn8SWFAq8M
bvM6j6WPZ90cqWZno09dlCLeT52w+b+zOOg0yQpEqZ2zhpQvTr1FIRA5yXpG2/82Ik9nagfZJDFC
/GlRfrH0S/2qtglA3NlaI1lx1s8hB2au3wDoJpY53HdGOwOibKdGGirvLf4MlT08kg1bo+A/75vl
QsbIqb5XpLYJ6AHGZQULxo0+e3uULwwDpqof99zaa/pQDvNm+/dcVqDFY6Em/S4/YHpc7C43kxxU
UHgTLAzJzjFGmaizBIu87tFy8UD5pMFxisEarlRaj6hRkF4BEIxI8qGgsVrJXluLXI5D2GX7nbKU
zf00Ai8aSuRfXrFTBNUIJQoDoTy2lMg8W8C/ZPAD4NBq/dyQVH9dNnkPx+wUjY1lK5H1OshHJIkD
+NCr8jbmYV/nKygQw2Gg+779SFqtYOjpbp0C5mASn85ZVwklwHv4Ea2PGoUiSWOT7yF9EwF+uMEy
lTmD4VWcaiZ8Pumf58bOPUkkyP2OS2yW0LYL2eB3GPDYADNF132Z9fD3fkh94nDaawV/QEsrFSQY
cEqqVTCKRfQwkJmIxjQAZ2YOEmdyajRtLsluOwcQvgwfYsk5vBrK9akyzjTcTgjloRqlVieP5bXW
M2EamgFH1zmSfeQW2lhHcERvNJONv13Wu51AMed7fUWInN8ULlrpYmxQOfe6l2ygfYUwGTztUnVo
5jrqfLrsfPBQjh957qia1TvXyFUJXmpAKM0tArFErA4AVGCDI8PhO9/wBldC9nct9ifc/Y4WNQ0v
DjHqEUjTEw6BkeVk1Jrgd94xNBkFP4W445lUYHpMvtGxHeu80xNtpEdHlS4aTLjibY/h7XhBr0Z/
kzPQRdVNHPzO3JKmUWxax5LD1MC+5G9FwLx7mGNddVqQ5F4z5QrPiZFzyoVJekAYw9XZDW4BXx3E
HU96I/a7przhpHMHdSMtxos1VR4FVMun5TDZP2GFXvpLVlAvsf7BIkn6RfYoZ6GFe8jfC22RnGz1
5cbj2J1H5YmwTE/d3zoW74nbuV/KIcbs8ud4Kglf5usG0QyTf/pzT79rbfyhjHQ9ZV+f7hJ1Toji
dqdAIFl7sNt3ReT2t4qrKDBeuitg8JANUEMn6lIJra3r1d7bsXEhuszw+y9WU9dDz1qJG/YTdPuq
qMzEzMZvJF8jk6TIaNHiaiUEWpngJBB5skmqAGduKzYyTCUST3N1mRh309aO46yYnm2S/7PWzPO7
WRAoVfm3vIQeR6treWOlRl8jYL5ZYZFP3w0Hu2uSAhyeSB0RZ6OG4drG+UrPkZM/RfYuIZamTAzd
/lASaya1gqUqk9A97J/dAeCPdRHGckfc3kO18KM2x8LTXauXAiBA0BHIx7hHrsFC7l6kn98S50l9
wvWNc2cutbWxRPRMxJXnANJ8uOxHA7SUd7TbX8FhjJ6gCsaaI0HK9UHMNyXAcEm9lqh/MrD0NyTI
RIgU5tIwC0QdrUcPCgnjdy7GV2W5tQ8htnFtFA/F0HJL0Qd9JUKk/4I9qrNaBWn4Z6ZqU74VpEPj
e3U3+n8tosI0DnmxTbY2TOR3r5HrhApminUZJZ91Whna96Hr+2q3hk0XGfTfdyMqyhS3Hh7BGiK6
MQqtcTCtDoDF7xqAmdPcF2ETCCd5B/vSKSHAJdE6NQMMl4vTUWHspUsfqrzENKOh5Veo+PJLa6xO
+tzmt04gzpRotRwpZ9iZ82iomg+defAvbNX0aOOqdRi0jz2qbysGBNB5W04Fa76/xI1L8uKFWiEh
H5+MH4J6Oo/OGqffPXrpzKbOSEeyj541r0ETUNgIR1Z2aiFLYJIJ/ChmlzJgRJFlnxsSKkHwAupw
wPvJdL+3N7la5VJtG/mIa5UWp9Pi3pIbHAhvEVpqygNFxnIjMZ0e39MgQLpVrS8qF3T8C1AohXwq
QO+d8xn5/P3RvFFuizCVqERq7qgnx17EQFAKPeDLmD/IT5GF/K8VRq4p7bDRjlTxzQB8QEsSJ44P
MnLzs2vb0+IQevPBdR3UjQymSmBILxCJ4r+XOPgcZtgeGd8qMJnd241GsX/fKcdeF2FkyLP45Kd3
8bfizen9CphLaJt4RAhHwZ5fQzTNFHMOH+HG9S/+xWwWW/SnauyBTaVXycTCJpONw6qcwwfgS8zy
tKzOBAEBJOOJPfO0hSwfUNR+jXbFs7vDGZR5ix0IfHAcSHUgxCtUmF4ruSIrbEFub/dHVJPwyVC3
dxh2POCZ/tXAqVpY2uafDxdDNx46VFZm8INrHB0siXojNBYd/TXur34kOa7cQ8mkmENeuewKC0wd
VdT39WNu/Hb/XqUUgXN76QIa340PhAVxiA3ue3s0N3PCfGK4Yq0bLtCEZ0Rl1wXeAfw/J3Nvdi4l
J8lvsh6cMad///DVkbXEQ+PIZuZ6X5Ng8+85slazl8bhGPbUb9qaOSMEpl5kCTA3jCWea1g8GdtI
hMC8lte+m7s/ZQ+7qTXG5keYYlMhPweKAClm6jB7LxE03uWqq8uT6EcgNYTeHFe5H3Fz96IFj5f1
VExlc5zotdYy2gfsLk9WqrjDxPccYmhVaVlch73RoI+J22ksmaqfBjWqz0AcYKE5g99deRF1c6+e
sFaQ+gchCwsDK0ceg8Bqrl+Y+7CnPNDzv///02mZY7/HfuANyBtQ9nedEHVwVb+LrQTXKuObSdsf
7LHvcgJ/HupWABtkUq1RQRdIbKazmtwe/+3rQMTnG7pw9I76y8H5wRYZIj7UpKjehuuZhF/59ilY
BJ3+0uIV9fKwKfgPqJVsD8G3cLkhTfuLV7j10Jgb0km5uR4gNMBHiaHsIZ2Gbk/JLGnZv4JP5IqS
Ey+pNWFS3CaHgG3RByGWKZ7uFlihLRT/akburi8AKp7i5WCXwYnLjAnLiq8oQAmMPm+SYKhxk1Ko
GnzjKqZ7DZsLfCOeeSX58ckEZd8v2JX1CjTeX/b5nTApHEQOTiS1bA83sKxfplsJzAWUaN7olYA+
QBEll3Ae2A85cHnotRT3QHxJRZk+GShrlpo4O1hfG47oVBzWJCXI7F/Tw7x+5WQpedi7FBfgd8+e
nrS5mrgegiBFlZclOwftELYC5xX2UF+sihMdSvbm/Wn99U/U7p15n6XWUvJsMbYVIJgpAottBjoo
GiCG2sDlU13H46aFpzt3aZnXEHg4IQl7GOk/QCGmeh3sLBkvhqhP8sVFj62b2Z44FmVivh8mI/US
6T23rPcatD5VKc7ONZdvzdDPbPqRN/lrYOUPRb9XEoAlkBypQ/I3lKjU85tq+gBbXUQ1cZh1h72j
S/eFZt7OAo3ksYV+joqHFyRQMMb4cpqT5c7ihmLBEO99HeVl64q5KfuUKkn2BvSy/G7k8T0hB5m9
BiONcQbm6t5Ja5JCPnBJKAAhKmkB+IKQUZ0fLfE1sFsIK4DjASx+pln2N/T9byHza4WBNPaATn8s
hQUAne7A8plrUGImfewqMzJrVxnX4KXeCe6HsGrS8n03hsZgFiYLMVgxCopJz6i06pxhN19mdt1p
Vzr3aWtIEMgKjygpeQhihZafhWn4kC3gNfHAZhUn3GXj98SsvGaWgmIJpkr4si+b1ST558d2YW0S
/rDhZM8iwv/Qbjg9JhC7o+7F/GwPf+vNOihqIJbWvzCcfDDQsimWoMKQwjY2hYIlEJogPjlojhOh
kLdRAImMiTbDN7rfh5STTCoA7zV+7J3Dh8T+NxpJAZhjCDqLTg2wlf8U1jI0H94b3ly1sYYSlZ1B
vikL0OUYu0kR/8tvmLpGYup3BTXZn/UUswzfEPql8lJC/79rL1WUKF3gljyPfIjA250oeSm+eJy7
aTasiqss7uV0H3Z002DRh7A6Fh9SuyxWxI5hdMGYdIn+vv1xlDxr7zEBuzd1pV31560TX/6IzRZg
92/+uf0f2oJl6QnC00+RCqKH3R62nPAfFRRtK1TSa13VYG4vElMU/NmmeQHfDMTl8mHHOYb0ZzOZ
TuIesC1Qwmma2wjzz4mOijld8Pv1SqStC3qxD4aY4nAi0Lkf2Wxba35wF+0VqXtZryIys79k9O9F
lwJ9MU3tIEnFU8XJ0RmEHY1OKu6t+890QMPVc994Dc7APEzFTR8C4z9OHyHOTadbKkeMFGohz6us
w1JL7igIZU7+JKvCcwoni+CE4pDDlXb5ut5VOa6SM5Nxs4J7i+lgScyGEMUJ3Q/0J1Aft6bAlni0
skxLoq2Ambyn4cgACCqfu/hiqHHdqVAbEmy7Kvpi9lSDjVb4MLnkcHRh0bEwTnQ2JN5rBa3QAVau
HfzQphzVljt0jvrFA06M/HK9rlIr0AKFU4YXGMd5vnLYvC1qb1ZWdPnHDNTDf4abwuOgMJxaPXyQ
6keh9sROxAYabxc1YEGx+tbJ9OMF0znjj5kBh+8f6BCVtTYmBW/UgYh2deQdZCBRt/J2JSXoc8XX
fNKRj999nIwXxkFTaw4GmI6TFSr9fxUVYmztFT/D8OCtVZJrRelaq1NPkvo1fWgYEA0zEqCNd0dk
R9Fa6t1mxesEq5t43+j5ukj29xxMx3qNmz4NXA8JFJvmIDEldfJ1GjtYfwUnviTqrT1/bEZjMKs6
Bel/nlqJaHYfwaeZpQexyr0TNW1lLlsYwlZ+7pb4xO6OeufTOPX5Ul0IXqTtQx7d+mk84kl1yBS2
3R9o4Ac32PYPRJDgLnJwPt5wuF/QXHu1iY0fZKL5gs5z6gZShT7ZUPlEaIfdPkwcxanZKm6V2sqh
PaMZnLVlRa1Sp60osT6YinmoWcwAOmh5+5GUGydvQE9k/mewjKFeQvptTwaWZ17knmJsLbPkxcx8
4p/HVICHB0AlrlHC2NFMBjeLMh5Tof7LGiD/DqOjAxFm/aNjajYLjLGU4vmRR4yn2xi5uiopB/aE
wtYAmJFv56K5QPVje8fXEP7fF/+UHsiGkhSh5pPTNQ9UyD/+FfdO0dOShCpSvBizyT7kfObtuilE
OT0A9bGOhNqgamlYpABbtWoWtgRsMRDlpG3LLUcwy5i/jtdqIqlXm4gr4peylPedF0HAPVz3PYS2
w10uwV/1ZDPNBkzVe4IAcnHe0dKR3jakWrdaZBftzrTOjv+gTnt4hPJSlF0qdp3/3bjTOM/LhwaV
xM6275LktnVKBBMDPwQwtM7BFCOwPATdx+m8OZqJAz0fFX9QJusbVYl6U282GW/nWIytR6nI1r0r
EuVWi6XB0ia/JIT9G6MDGCqHaa3QLjFXH/nsHdyX/SAygjhta0/JBnAF0yyVhGXN5xpwFUJwos6u
J4K0fjkZfc3NP1jro7kW2AEyqQbEaLktODtqT0e1/Q/kSYOkAqetnNo8d9lvXBijKxJruxUFS/47
HMtv15PGeQ1haJTZuUXbQAdgr2yhwGOsGfwfVDvbL5o4QDfSa9ONhmJ9g1LyGudnWhCCOVKMQVXd
5UKwBPeGUcCeXi2s40bJH+ggVF2ZGBDEAbRUoBsnHF7qQIbyWjbnQS9gUWHv2B81MMJRgjOVhlZO
Bic6+rb5EleYRen8KgxttIPiQPjMm2d9BsmRbLo/08zEHTdfcq+hrk0HbYLz5zmVlDNv01x2H9O1
0+V1UhIOQCQRyNoBkq2zysMJKjUzspjjQgw11TdyA4sd70JYkzSnzJtxeEtmWK0N4hkqmEXzkejC
hwO0qG9Cuqq2xLqlAhYzqle9roOUChMVAmK5KxiI+PT7D1wKezkTZTNzIZGqDn125xCHhRiX9gQu
Wn2EijtixnegP6cwyu+NeLSBUF4CaZY/kENQsSjwnHEmDStK20dwKWEQBCll3OI26ijQ3G0ha2iG
dVYRhAJrcUn+DuvQrV36rx95/uxlWPrKcsej595pUF3MD1qMtMl5sYpUsRf1vL71Tzgh2Qn1aMy8
9y9NiqVAmQM+lyrjIqxi/InOFKFMwwM1fFB38re5ZWOoNes6IuP6xKb/VCklNk1nfO/hggrWd+/I
Xinf4gFk3DuJXYWmCrgh2zcF20a0eG8sDAmHcUjHc8kFW6IZ++Po9HOpXArqa7xC+eizHzzVZOYE
uFY2b+1eh/g1YrM3dowJtijo8YUmFRsET7F9owGyA+PFfjjXQ2iGeTWefYdMXg/X344axG9Qipxh
+OAjUosfArW71ohTZfSQmcoATOdqSETOHqPMkLGgRGnV3+uB3tFzY1/vJry0obyqJumhcuV96uZS
dmL7AhCXMZFjxDgLglZBN5kE91pmk/XAlTrE56mU+RCkNqTk/l9Fs/M0gVYqrSopl+RT6rL+Jr+h
0FeCepKO+vzIwGv+ZxRuRhU9SdUDlShIvvTGkGvJ0VNZGokZ2Q8U4I1+NihfFppoTKhTOzcUnLFZ
OjLTmCfoL2e52jA5N4gfCWNT40FiTV+5DpxJA/K5ABs22CEhx2Yka7nYtNpLRtcEG0ZK249kO7NR
UMtEqKunjEqFtgdaTbQrr0Y56xgsHTOrJQTHmD4rXjlwv6HiLuFHgtdp4M+PXYPIzxt69ZVc92gT
5cgqH0zBLtZo2z1GwblgylCp/FjT5kOg0HzItxqLcqNhZr0+PePNMcwIU3uvrmHCpxbgU7sf6qM4
5Zwlk0n95y8c8kaC7gqGOImV2bVzAYX7N3jLcoLg3pE/rzoIuQKZ6Eg/cgAss0m4LIjrLTLNcsZW
aiUfc8tmQrxgDKq3nSr5BvQSkUDQZwuF+6S9Pnxgp8iV8HHITHKLLMAEv04QFzC9ieiGs31iqjaJ
GFh7l9yeScblqOA5xltYepncLzIU5/0a0VS5uzRHr0DpeakOdp3Z85BpZjB3+mhROg/eAUzOhupl
6PWDJxWEUOa5ZixyMOhyG8gUaQ4soj+9mOGw5N4rtuAle/bk8lCCfEHf9Wf92m7aBc75EXsiN+6L
QTQf2iopTI860EQu0wpqd6NnZr+vFv9Q1Z6ch2tAqkczN68XegsxrNXzRQwWT+f5vRZ5IPeQnKKs
8xxk6TLbTELzgZXVVFZts3ar+PNMmDopeHVV6M6Os/BB47W77m/X0iFe437DOvLMYvavIkMqQF4y
YU8UkLsQXiZTKOYsjOu1a128dWlit8fNn1hIPa0qiJvHhHG3Ufc4gESmAP49+EP4O7TD5OmlEyWX
HNyeE/fuzHptfx2n81xhFwYf77CseYBoIy9URsJZuYZeS92Go04XRrAyqkUMFC0pYaKojvBnORJg
gz1BuHJ5KnaQrc42pgJfG6FLzFPgShL6k3aFhFR6MyPK9ilxOqaUcWy4LaqthOxwkKJl/jbjKu0j
keGpnur2gqbKoIp0Gc3QaKLTe8vhFM1sgx1VyYezakxnfYnc3o99VTRhH5oJ+1RMig8bIh1vP3yn
ETXZGiQnees7W8LCKPBhm37GTtcT4vvVXnPcCDFR4IrgQ3L1ljNJ9GiPyusmqmwFbRZ6Szpv/lM2
WTQBQW1WwhDg0r7iZE4AdQNUss247rhamu7l3i45sYoDon4MNIPjEC/x5mtM80c39T0lz2BxJduy
JDVSlJSkqZyfvSLN00LTJxyAmdkaoMQZwq3QpHgD/vqxlfQ5GVnJToJ5ZmeZ/brNaV2KHdBCs5yp
5TFS70rdLyExlYoS4KtdI5mM6cSLCbl6NbuwkakYUIwYHQOVdbCbcicQGJcyrZwmtdILZ5Mb09Dv
Z9RFc9UBW7AHzl0yyT7opSDxowpXaRC1obzSo3X17OZvl1WRJPn6iJuRVDcXUzwOAcDh+Xqe/CqO
CbKbrva9AJNvGqbkDy5uIHqwfZYuD4nNw9oc3ASOkugJJsbjdh7buWnGxJo2cfjGmbORQj0Qs6NN
AYNsJUkLfmXHDFC/gf+8rC4InHYdiQxJNHsbegtOTnQ/cw5IJCbI0QlWTxiz5+7zKm6ZIDuhBqO4
3tp5yhupR1PiQ1D25oSf7R6LIrqyHk5N9JMumYoZrA3vEE2uTOQJWC07MJ/nW4itYGTwHtlDLiNt
jBnFWBJpqLVthb+t/IGmlWYb9r6x5lHlxyTptfPknCnDywCJoHtTEs5qfJUVOaNlYrsQJcLvCbsm
KToQBFTy/saHMtP77IGwJa+dfwNsF/vYV+7TlmhKkzR5MVrnztOQRIkTJZx4Q6bwyzwRKW8O/39V
DXlXUbaRlO0TK2DL/+Kgc8V08q4q9CmzP3hkQ1/1h9nwtOs65q6R6OM/P1yqO/DxvnZFwLjSq1sL
zOwLQC66YfyACWO2uHwPFXKNGzNzti0Nt7v+0mI6RzxehLz1jdUpuffl83gqtMO00TTfqbDZHNrb
HxkbrQ+R8EfgPKEJAftnSygJO5m6TQ5STHt18jJ/w0SOUlRUmOaEyxgF4y8JlFS87xG/mZogO+W0
arAxSk2LyhpEo/ek17pEEdoUCRD/HckqeXPRaQzC/31zXeIq0jT2ZDg64hsYtF2FeC+p/wt3FwTQ
VQbGTDm4E59pyhfSfc4pBc/Zl92g4jRJlbb5Ko18PfPrA4KVfvIZ5kiVdVEvksRffPoaSpPrlmb2
M8uz20JKZM8psarqLfEDw07xnvqeI0KeRYDnWvt53FVFs9On9WpjYcqHea5qeNfemvbisZzXheIk
c1Nm9ZsPOV177iQypDZJTzgZPX9+iajGohOzmqQCMoNsQFM/GSCvwo8Z21S+GU32gS/W0NLMNS1N
Ul59ETdsRdml6+52n1wpaDGmvy8RKwGawngqN4R7LGsKJEhSwUmRqIKumordtWrn8gNhgKkzaTKJ
Rp4mNJhftNBwv39x5vS37Cen9nXnUHXmT8A9iZoX1kzOC95ov+id3Ggdp67RxvLt4iC2JanMOPIl
aZSzb1vCoY+Xy7/uyZemxWuW7RP9gdMvOuQfAascibWL5EowUUfVBOZHYlVlXoN0KMCyv2O82jpu
ZBLD4xNsO7PVFKJf44HVrT1Ld4d/bj4IE3nM0e4iDQjO4mmpvWDG8rp5xYpRlB1quL2oDOLFoS+A
JZwF1HhsfQO+zUEz8c0qyKmdoORuphocGwS1clGj8fOa41SZtLKD8ZCZ1W9PiQmo4srymwgJfW95
LwRnhawbBj4JbMFUGGKYQ/MS5QZQMbyoXt53txZtki3kEVXMFOyi6d6M74uPO6UEPKWDqVJ4lR32
1w1Ivun8DegI2I9lrYQw6yGOfb3u/WjUyxWDuP3RbevFRpDbqQ+Y8gKRNntdrsEu0cv8iuP6x8Id
JNo7yHy8kGaqvizLVcyCAf8znU5Cj4Ktnz6O2eJRmmm29B0NrBH/NTOPPDBA4jxzjSxgjBsV2iYX
pdFajOybclLwi0mNeepJl5bmtHCQgBwdy225IvXu3icj6hFmh7S/YIC0yM/naODVKDrjTeOxeB6F
y06W74ZJ6qT0ppHU6oemp2fYeqzZM6N0r3xs5dMNEJBLYKX7vuLVkcVno+6CIvxRHCb5eMdMNa43
dOsOda9dTYmsDNEtZI7wuCVBRVwUlskxEJFM5HqMemfxfvtRaWHSlC1yXKBP3JYD2kJwtz7JWsAs
siNTf+Dqq36/6+978Qw32UomTZS1JXaPlYQeEVClKbfOz0Bf5JJvHjc8RqavfvA7maW1rR8EVGIW
i3ELq4d7SMiUrr29Vqrd79dwU3G4Un7ODYqpodAAqcA7RA8cR8o0FDG273QYddXuQroeHoePiUhi
XJOq417m3il59mq3gcbAgV3OPgwMov24SRNlhvR9j3AMF0YCfFcq7gnMRGdJSqbUsiFEMlOZgYiu
dF//qIudLpocNl5LwqPasofUiTQ2FjM5xXxDKwH5C7xKyEAImuJYxpzffZ6h2d9SBJtKCzt9xSu5
4dFVYHx2etvbxbU4CwTxb8r6zBz+cUXFDWFnI3etYK6YffpmXKKRpMiT/NwoAOPVXSpt2FEWCUjk
wU4HZc2lnOaIQHu1LiQQqpu0QGiuVoDlWNZ1H84bNwqYE2obDGpKKV6QRnf+hOj9URav9bX7VZIL
620Ww/k54CybNSVw4AGqdMIf4sCD9MQJ6vUdVji9tFDahswWXKEzeCDaVZ34gdVVf7sx8MJ6XNfQ
onu+gVT4oR2VMWOL2ApKfDLYolQfzDs5sXuYFsop6VG/LeIkqj8AVAW1MaW6NY7QGaotWBqsCFQs
pPSdxghwxAjmR1p2zXBSOgwPdXQsUqedcQbRNZk4Nd42GSLHIcZiNO6jQSNu50ABKoRK+rexxxmg
ptoIzN9+0M15ZRZFPviqYte0+bw/sG/15Q1kjNMv/PvoiJr+x2Tg7EdH+U78B4FMu32qY9ZplWaC
Aet7G4amRH/zM0+QH48wTiFWMw1H1lJG/mXJ5BeLWSdF60DFu7iduHmPcheOBRld/m/Qm3jOwipg
AZH0TztjuzRUGUpB/f0sTAL+wuoL4gL6JynGzxu8XQ8TJxoi7xyDRmTG0aSBQZGVXE5HkQonwJJt
k78w54gh8wVfj/G4j+J9OiJBx1Qez5jzWFpZB6N5Hg6auica7yG2tdgRU/uH7H63/nj0NOx9C1FP
uaQeYfATnduOpWeLkOZJlIi0RhcCgUfpt32aReFFR3VbWUcQoMdBEkGoqVC2nk9/3HSUhCUivKi1
mAbcFL/512agc7NrdHcDy+dfHoPN/t5RYbrilg7uHJKeSDAcEgoAVbqduIj5uNNzt/paWs5t60ec
tz5mBjUHJQsBv95k9D9hjEIzNuWmnDtoAq+mnWqslI7OFpTLIq5VDIOYoxTzLjRav30HJmIyDjCa
IHpXDoFD8GL7TUNSuIKIm68Rob+VnzQK5CWitgwmue5kp5QTgYigmMreXXorOQyrKqDNGisYwSIY
FCpk5XwgpqSmlE0CdOrF3iYagNjr6YzZhveRyGOI+JvKLizHy5L4u9SuPoVWVlgESLvHhOhu0La3
YTG7McbJCUR1csfFzIeK5MTqLOQcqzXMAU/NyG6f7stWQxXFc0nZQExTJB8wGOIgqef6O6BJu+Pi
oQKGfAfRAAzACutnwE5lnWlnSFJUF1Bx7AK6UBnwYk9BGAM+mhXM67twCTgGE6LDxBiUDqlsdOoN
t64ZIjOT3gNIe+l8Jb9BnXUV6+Q1MbhmNT6JmecTuPGcJugMwMecI1GlywX8AqNZIpqtsOnS/uJR
ExDcd/rBQX4JbyIL+ppRmeCfgHzVt/tINJMAPC2HYaMQHDpeDXpnC9o4RGTJhJoBpWSWZ5nejnXC
cNf4/Bz/9sE/EUiQGJ+BxOnRwpj6I4lkg6qLDpq3HniiAfNV2VjAhUwj44MKLXkgA7nY5DwOPiDK
hQKn0eSCh5yHSbaARdyd+QC8Lr+78gUTFZVggJSZzAI9eEXKKummBATC1YZbPDfnfnGTq5/JqvHU
x0XR8ysFiOxRJ9u1bCYDo8FIh4PI61SO1N0aOTNy1LpCbfJUT7Om4NJP3Kcag0OBGZJCQcoNaATg
VdHFY2XUuiPHK0VWFyQvZX7iAg6d/KpKy41V4zmKTha2QSkDh2XU3Em7L5tHNi5YUe17qTkAl/Tx
6Z+wVZRjJ2ZgPrkbEjO7l95fcseAeGDq3nOlLn6cwrIwRzYp0cJlA+jORnxwYMPRiVspzZcVAnGi
EQzch/P4kK7txErvh2lCT3YTBTepuwyHLB38tnsoydMtkqYSWwJ0KWzU1P3bDeTUa/PrLyMn8sNL
GqOiG5UbPvY/sdCqVq3B0RNNi6KSjLcPhWvV2GkOw/LuhyH49F+pI8tQ5eyCkYYEyTJnFyqXa4qQ
4SqOLRJlzITyF6ABXTa7o4JJzzdKfXCYzFmwOXo2FALH7gKcWy4qAwM8kVMIh1yrXKaWwxmBTcRx
h8qkkLAj3eWIT0Ah2u2P0wfpA7MAv35K9NQDu/4vpC6qYx0ouhLLDQuG/jZzwwybEzjOWIq2eK1/
oC2C09UKEYhcdKLAnL+REyW0xdhOJCbhGBthqsL9GXSHO/FwPtQ7fNKkA0eBxmAiw2WXWm65GvZR
TJ0G19X9xcIuB8Dq6ZgDAE59hZSnfRThJ0nWMcEkzOm3Z6O5o2ajThsuDD6D4ycgCPDSpU3x/Ba6
hRMwwnDzzCBVkXB9ZY1JZzUdbBh3P8oM0jYqrbocuv5lTVzpVEMWygBd1Iuy/F8LyM1TU6HnuTND
VgyUAqmhrqpxXrP0ZPR8NHCRvmI+QxrZ1T7d7g0WN89OcnP3mou58iZbdOFTZIq2VLuY0UEtRzEu
UntpYLlYNUMaGNFRLWi7Xss1VEjTx14xYtWb0uaLC9M1Meo9XdvKh+gJ2aU4eaqATlgcubPntJih
sWuqjMFE5v/8x65vI0R1si1DwzJps3FbV4XXMlJ2CvBVciPlyOmw/gcA5JoejRZXQ5ePED9ZXClS
KxHkpj6bNZ5TKZ7CbP8qzAraBWjHv/DFyBTAia1SM0YYzSRtcNojlyObfRgdT6soGsC/lAxknndS
AV1BA+pAjeYNqa2FomR0nRp/g5d5xiz6dXW0c7juVRu3kqjNfffEGKbR58NUAkBmCStznXzi3xb5
8ALM0A+C0VbE05ax7659bJIci+mzSGOQF96+h+ckZxVUCJ0PeRgngAaXWT8kKTLuKEEGr9tdbcug
UI8pV90f0jf6GS0OO/3y6794S0Qk8Iih7nRchAaarnjKlfQXq2BwAa9dt9MbYVjvSdsPo5O1sqvk
caB15gl0qv7VK2dVx0bC2c6MlDUsEEHCWnLiP93qfG1lnMpJC676kDDy8nYs86S5GPU92l4xRmiN
HtvKZtLTDCWkpkObFBBT1njeoZP0zc6V4cnQgqy3YXhSA345Oc3yiZKkjxRnbVNAKMU844fbSIi3
xgqkBoXJP2W7vynkAqAJpRn6oXOoh7EGT3ZRl9XNWMlctyv/3XtmPjAyLpIDI/BaYn5I5b/VakHk
ECBhGXpBP44iB8witeyraxhHzv36OGT0OLIGdDUU5gr8fLbI7ajlD4fhWauAZPMyK04lB2TdGlAG
Gs1M2CopVWHSI5ONlpYidH+aGNDOm9FDcgDvm4JxZDbX9nTm1FLPnyOIy/6p7EmFB46u5KZ8QNoP
B0E679V/+n9R2ksqP5f2/TJVGNTbXoGf9j9JT2zMiiFT0CLwY5m7SoRUt+VKrR/KIUyQeS14eegM
WZI11daWRRcq6egtaN7j0eZZIfscqwuQbjAmJJvnYaZ7pDs6cxMhGdUD5rtOmFjG9HNqMs0GdhmY
0ZSZVAWC+oIci0Rx+VXiFeywxAPQnTeM3s7zOot4tCObDEwuKziAYo1mk1yOToakkwZ0hSN+TeQe
y+qGWavf2RCK0111XHRwFUxILPaIXUCRdtWUwM0i10MEXdUzpKG2QmOCKtz0MiE8t6G0mNZHyLMF
PQ22s0D6Z5PfkhRsHoSeUKZFDlD2SKnz29prXYoc1/ilp2a1z4GB2m8acJKqN82z4oK3lw23uPxH
oMpecliF/zPL/iPenhGoVhTZhQ4gLEO/R1pf6E2ha7nCjNQmMOfd9p7V7tfxv4TelHzrpN+OjhGY
GLG3yo0NLqaCLkOW2HDzFhhB+dDWyB8ciaZNs9v3jec780Z+ciCTS1tj36OR27jAwc1LCf/UHyjB
NTxNeKRjYUHHV9hWfes6ArQLxwdmotbajfuYifBq7zNP/z9+5rI1yimolfoqDqdtYeKlx4tO+C3u
WUAfdxZ6aoF3sGLpLK4r7yLyqIEJEGTYuMvayIOLSHi+5At4f2Ok7UFz4ZDxeDRzywM8cRXVZTsW
sVUDMMyx/Zor4FVHLV+Gos1u0YynuJ7yBw1phCFkMSb4rMeXvIzHA7sq5wxsMdJDfn9ldfZdog7F
mlvPhWFsAqHw8MbvduSWpPNaPzxTKQq6j7i3vjU5iXYg2Xtb/vxHa5HG2gZsnZ0omdnEHz86bTW8
Eu5HIyjexXIpBzicOeIvqy5UmHKZr+PmNAVPj4FVibl61oNnamoEGEuKjWid27B+a1i5+iUMhvYb
ulntZtj2rHfe3ciQPmV6MO5zgeGaT2Cjorx46Z9BJEqWu25CUgG/IntpM8WMitDUruMec078M88Z
JoeZXlos6s74PMWlsnC8L1xq7ftID6EdD9q3KOZCV+KJlQ407uRD8oL0ZYvYlsl2LhNp7W+6nkGv
m4RtNxKS/9UQWg5gmE3b6Xl0B16ccpSnqWj3fgDzWr8sMHKtdp7AxFtaRyxC8mO7gPMMDHZxe75a
8QMMk6m/FbOb5P6RvNGY5caZ6RbLCtS5CKIL62W35DKuttarI/Zi498Ut6VDX3a9QKftgYFxfBhK
IOn2smeAasOKt1G3Lh0+f7uRjAB54Ef3G0WGq+6+cQtDlnY1JP0dcS9WErSxiuaLWveB7sYz9DWS
u1PNbgRGOR1fpJSvabImzLXkVYMP5pLrg6PtPVHye2V4pmGwhN0xjjsZmow7tdGU/wwQXv3egMx3
zzVxbEQwfDEtWn7SGxCmZFD40y97VCR/mPRjpiS6AcjkZZpytYmCRkiGvpWemAis/dRyGF3qvErw
SsqRv83FSfrLEKGJye9FABK7UO9rgG0E4vCRmr+rBd6QaJonXUsQqAujEffIA9ZwIC0W6FfQ1f9Z
pyiaH1UZWxPGzQccf8tZnd+mLCF4SS7D6QtX3Y+A+QIUbnNeMj6RlNwurwKuexExdEGqkDIWfbDl
0ckiXQoJN/5lPp8NmyDIshyrd44gBLvJGFfDJSPrQLhGNmNeIw74hvxrKpYsaqnMUR6rlG0Xuxcd
UgMOs6TjcbyRILUeaP6Fnrmb4g0+xd2R1yswxy1zUQJc6INZj/ySiYiRrtgnYyxyt+9O2tJY688p
/WOtQY47RQ/y+Fyjwr5ec9O52+awzPj6U7fxf0V76dULCht+OMVONgoLU1h8XyrGI/a6zghfq3Ti
J2yvea+c6XW57Z/mSnUOJNBC4q14szWn6rWGURpGTGJ4Ku0PEX+q1Q4FCuk+s+zCdBCcSZjL1+V9
GZ2bjE3tCAm10cErbbRtiHPoAO4nV5f9xaqOvH8iqJdXmuTji81fOoFgqXysRwAyolprO7oc73vI
Oc++ZKAOnbZYi2wGSpVDDldp+p2opeFn5WmmG/mY9PBly1kM10PhJwjVu8v9nrr6yPC7OQR+z9Lc
7bsIsUFdu8xIobsZyumMkm0sfgQliayHdFdHrJTe3qwz4H+/uE+ICCbtK3RczkrB2rsp2bWSodY/
csyhBgWST1DfLbzaEFbVB1M8qAKVJCPzzPnwTJjaeNA36r8b1IJuw4EjNffiMOhb3AmnzeTu9t47
zE9VVJbX3pIJwI03XOs49LTIGWhrGMzb13t+h5EEQNXuU67akCbOxJN3zxm6WoEx1cMURoF32Fo5
pzo56PPLIWPymLtTsAFKMc8YkA0gdOLDoT5R4sW7jrIZEBE2IbaI0KHMe23ltUos7YUJq43a8GvG
1n+TOxRgLGLpCSGt7ANIOgN7Z6LiShCFyv7c/7J33fWJJywPQ66TxqHHZUj8dazg241ETsuvMrPQ
l+OoKeU4RI+7HAqwayc1he8KU8X6GPrUxbdjFI7iOh41REECQBoI7eiPEx8+0ZjncZ7cfdIRNGDX
LRG+rn3wJSz0cQIAhLHW/0F7FC34U34XayyKvzjMpp3PrSEGcP4p7GxPcg5Z8NIaht4dhvLczjji
aBCdesHMvDoRJk/eAd1MeXIlHlen2z6b1FCwacu7LI+YN7ow66+rvPwbRbYi9kmxXxN88uoMt9uC
eiZoRZBzxYBqlGZYnC9R8OkMd84kIHelnfpLz8tIXuuBrRPAzlLMMrZXmWjHu6ITLp/3eRdOuFgt
X1ooJ2uuUgUd28PgUQNV50momTK3dIgnwY5z683hGPR6k+u+K8uN5tQPe1aLcZN3Hb9fiU8FLAuD
zeLy1zKmFj9vP+DvCDvuD7BE5+9474OxJMZIZKzQI0XuutIayOBF/FYGP6oXJEgZ7fpV1jvX+/oU
AdsppcqbZh5JBpLlmjXJC+91y9zSNO2SWxfyNEnCqUiLYV+OVHMDedpLnwJXO5j2Efj2z88PfnxM
cjadSZPo7EkbfnWQSzaCzD6cqH8WpPBkrDnXsyEJIMjxzcbDSD0Tt4rYLnaAQRXO84pmyRRra5fR
lf6nxkS7Jd/4G83k4CGdqE7fU9oeo+zZXnHZ1tHGzDSrj2VZ6T6UTb5TsXSp8AhukZDfjU7V9PTU
2FIOaGLVIXSKp/QfmRU5rrUPPr1rP/92qlqXJCUQ8tp9+bYRH9Ah+RBAmyPKC9IWSdYqjdb0RtHq
Q421zfqUloE0eSIz1GtcYCH9g07euHkXuJkY0BjDBw00LGwie11VALjIez2ZGZOnH1cdhs4Fz1ih
QDDmgd9VDkzm+171l1X1LFOmFg3t2Vq9O4NLavOKkzlTsqn+AEPIn/UngW5KeLa6zZaOY/547BGq
J8iQFIxpRiRHE2Ycf3JRIPUe97GHHe+QR7Z/nxEE3H5uPHKcXog8NmxbX0mWmhAP4JoNYjiBqzXy
xenD9bZbqOolNbzlVbx3YDDmiz35+d1Xd+V/s7VHGvUmsFo09n/Z4Zoog0/+GOgS+m3Q25VDPQmT
I+FHP2SWAOpmhatcbpvXGw4tSrd9J3f80+P363vAe/D47ixhECXfo6wgIk6cEs+DkqMnqk3nCzMB
Omp9myyKgGxlIJQqmHlGfVUclfLKpKlVKj1bP3XVktAVANZBanIJ/PowdzpytZl4LOBXMhc0Tg/8
eAeggpBi5K0ThCR/LXV5OuVR8/NFLkuHj9WzDo9wlrT/sgetnfLkHs/R+HoD4vmHLW5qkCc5NyFu
8zaWlogj7gqFDYgeMl8ondBIiBdnggpA9Zla2qqmN6P3JcnmHKfL6tKiJLFlWMCTL3Ks2/4FM+HR
0/leIuCxs/bsr+FoYy80gn3POqshTOYKMenTNURXAhC4G5OpRfRTyTPYsWIRcE51UOA2f1HOVKDY
QiZO4PCcZcrZPzSW18Dx9GNq6800H9imyLPTIAHps25k1lWuQCuAA0erarqf1ymnlVc9dlgRjN41
oatnDB1hwtBfVKUKUWNRxRATjAaV/zC+OOf0WOSrUgbkyu+bP9ujBR3ckPmsbROT/74fuHfXLD7u
k8YuB50Pub96lRMSxjkZo84yyMoBB6B/rs9JgLDHn4HjWbgksvRS5FHEfBXyS6pPwNkSTi2yQBOg
2hlQ3InZQ+48ZhshLkd1S2PoNh3HRELUted/vrWfJ5VFqaUXDFzGEbxK/LVPk0K+RNFmEDNf1WvZ
OSOsGK+qmhlAfn0/FLB4yYnx3GBQbsSrJKFXdT9rNzqiZqEMcyTCnO5u5SC0ETc1/aUbwi2JhHC9
iD67xRIW5IcXWVxOmU44/X3OikLqmY1jJxUOmWcABgEN+lVvDWdRQfJsC/TrPt9nH50F0TSwB75H
RsxNyxhi4aBPiChEwktWpfO161FdnY/fCaPIZjfsomRoYvdpmHspezIFi6smwyuL0IXtoVsoLrcB
dfFp92J2kDCWygdtdJ6jZeEebUyXv6sqayMS1G2/k+UJoVWL3Da1qrlH6E5AT/JD5N7/jqNEHt3s
5yrxi62PI3Ph0hQ8OKIVzZUEEcGDoXhf9cAaXStDzQyTHuEtOw+kNiYITI5awZJL1TOwjOQXnZl8
0sWzef0nVHAqik4Jb92flbr4aI5xRmJ7avt8/s9sLiqRvk1Au5Ctvy0se4lF33dWG2wT3WpN+gCA
3BLcEA2b5xpj+oBeiCbEH7ove7ZgvwZiF3YPLteUKCe4lysk/q3kmpfc3+1bHVnf5UtkxUtvhRui
pIA9QYZ+TI6gsd3cNjgLkxA+mrJVg/1OqrbGtG3sbgTVmbN1tey0Y+/2jvzbkHtUQU2JVazVtAhU
HZMUhccdJ/lGdS6K5SIAIWQaVnEpotyqODUH8vtl/1fZ7cdQLw4hjuh+0Rw6/cmxgamzG+hZHDvH
3dcuYGu/Cl/h21PGtjkkFqYVBEc+2PgOVdCniwfrV8SBE0iyvhQ0A69XwerCotCPj2PfcRb2RYN1
mP/nTewbjPEdOhAr2Svm8X9iOF3454MHvp1RmsrryFKVJsxg+nTI4guhZzkw6sTGX27ZrskzaaSJ
TUKFigt7vDhaT/zVSnGfF578qzh9Go4zABHnpJWxn7IAlN2KbzO2c/2Vbevz2pf8O6bYPyF7ZImZ
Zqj+GeoXIf0gFMEXYlLovniADH4gWwp7OzA3xzYTAZfJQ6kSiW2j3BuoC9NQtsq0aVjWmVn71tet
AafUCBZTtHQ07Pxze2FPxQ13E8vhGWyxDbRimpTI4jvDAM9wvLdOnYFPjzD9C6yi+DxU8GdR93NR
nUTpo7Qx8Jel+SZuNZp5s7Jnvyg4U1cmm2rveD7H81KK/FUsbeTGA6ZCZGVvDrq5q25ah2vjDCCm
1/ZTJ98VskjwqDSNgSFI3ihpRZLXssR/C24WwZeq6XpUdq1Cs/x9OI5k+NtM01sdeWqK+WTbL7ht
brWV8HtugrkDsF679pkJ3jYpS8ffgyG4HDFTClhlIryaMOKAWsPUKb+3V474ZlodojfCdCCi/y+g
j0YqzANZSGe46ndSkmBqLbPH599TLfh2Ts9aZwiRUN26tAUbqlnSNd0nUZf8oUsjnJFGahOuW04v
YWEnoxb3GZrSJGMa0JqK2uubiIS8E+n+wrq5OdMeY5HjkogqnyVSp1SmYgN5tC0XkS/eCWge1ImE
p52hakfqHq0s6P0k8XvRGLysV7CM2ujVtn3hXqUjcDtGu1jL1Fg4X52mqk8mb1/Qg5zX4JDZLSRq
DmWMqQxOCToocZYx2BycXuHBdqpkyG7KPAVnYciG9marL3Z+6gxZ6Hrhh9O6G0irQYKkrmPKg1+u
a7kk+fAMe62qgRMNQEqv17kYIE7pEP+cQ7R9wletc+9ISMPcPTok8OJxJpMXQrnpwIt2eYJusrHu
RaTY1idAsZ7upoMqX5v6chqzONPbc40hi9BkQfSQWT+zWcM7EuO5YSCUIlvxt1z3XszS5/Y9XOOB
NpW1E+NdLu0I3hg10ZMoISLyzE4YG/VKcrdrGzudaxkIEAMQrOOdy3VWL5Lw9OnbWz+sWEIg1nVD
cSX9f6uht/WWEYcrcbxXiG2JV2ST+vrIvhNvSFtc6Ec7S5s4GkQlF6TnXReSm6PZs4a6ooyd0zIH
cwSnfNVKg7f43b3vPVmVvoS8TQpw3H3ilBDAVT9Y/jfoHFzalwuHfk5oQtNivUZsMfFcyJOWO/lq
HDQbbFrwmYtYfX27zg8MbGtOKF6Vl8NxHULX/RAXfczTv7awbagVyp6ETiXOA+bO6puOHaZ219TB
pYiIJJ4DnegsHnYhQiR27lEalit5qZC4pdUbBJfBBr4u3Iv1rblJNJ1VAgHcch9a43aVyCeBpWK4
6IL6KdEQ+rzkqY38ZuNOg+h8eF9mnw06KCSTvc+3qyZBrnVWGnAQ0KE1+cUs/E3hVDdlh4fYuBIE
KhwgZFYUq1L0bWskdO+HPQgl133Pxj1eksvencCQ8ODQ8gjcOYnNo6kjI/+a/Upfm5m0J57Am+ol
OurppOJrv20glbQZarSk7DRUdkjM3i/KgIQKk/6cK3ZiOg60nB3TTXd4Ddw2O0b6ep1ycYqCaDen
RW7aStcuvV2xhhjmAhW5WcZfNq2aVfnnT5ClLfhrZ27X14rGigdj24PEYo89z6mcrJ7D17aVh09O
wNFMcFdaJ0XTzMZVJMCWmqUprvu5Ug5HNslY3TSIwOlU7cZOOgzV63Fe74I4eVYH2hg1AkMyeGMx
x+//87fIi1+qhhs4qj0nWYfj0eZE+lGJHAU3bvWw9zSnE6w5Kn8fwjboypTYakcCuS7j7hAnrSu0
STVWnYRKCuVfVadN46omRhEF3rfIMek4YZiVYQ9/QxvvdSBe8XN6k7vOggiAryvPCnQsP8onTR5r
2Afnl1UPyvwVTu4AxiyH3FWKHieSBolNs4CkvS87YIzMSC5AnF8UDzydWUiLxqGErJeG4G7CeZiA
nGTl20VlsPSYYuCgZS+8elcIpPUwbWdcx7A4PTLIwq5XdygER07jWoYsqtoZW5mfV5PWDf7oIguA
Xczm03zbbDdI8iwtozpb5Ae9VtZ4slQblnPX6wFZ1o689Sz9xwjMBMDg2j++XdXEU8hDXXAf3KRF
+e2qOkUKiawC8AQbcL6ETgtjHiapzWfa0PCCUx1twy0Ksj9V/qVTwbjalohkQZTbOb0mhX5etVE+
vvlaFv907jg+ga4il/v/qqbrxvbfq3zL0zkP6cUPd2opAqB1Ep33rFyukVz1znL7J+/abJM0WY49
7sA/mFEgQ2UEcHitMyM1oBoKcl7UV4R9bVr9kUyyig1wzNSDKRqrSSSrtifVu4vI5Za1Ersq+W7c
vSuDDwoCnVaiX4dWt+2NKfkEeNa4YAhcS6VaRstlOIqlP1O5+KvO75HH481nhrwYo1KScgt3XokS
hpDTnFwaV4fWmPMM1s5DIjL5Qfd7VFziHpCELCJybDn/e4O5hR9DWvO+ft2jG/Xb+dPBRHLHSfuu
MDkL/1/besF/CluoxtS22j3Td26nToRNoVIwfdKpx0qgM3CHdZlA9m8ZqPvCYrTEB4lAHksEv8z/
Ms6VVvzb3CQS7fo+yfrAvs2SnHNnI56UgY85+vxp7cmEuwwLz1knE3yV2Gywfmbd9VXhYiFFjur0
bgSYMMfStt8EqjUtUJr4lqTAxkDKDsOL4EHUGABj9Z2SIh5ygzIkSiy14Je6mJLx+dj7o5yM4KGF
z2MSHaJYkE3nPOiRZVDsvi9gONeWKtaKyxR9I4AXPxTpi1oVSujS41YllqtQbrQqcPI4D4+CBISs
SBFJ9KrnZMXkTdeHiltFmcm6cRkzyMCJpPmv4WzKMUOdqAeKXavC7XUpJqJF8d9Eaufl5wL8GBXz
x2KrV6u5LLva7DuqTFuOBg1LhTWANuYestY+L4ocydVNyrR7wG/IKzh+caFgo/RZDUp+rUKZsKHf
HodmDluRjmXtsnLWFTnmzbvW7jrZnHpktJkxE3kUSeqWXJNWkwKBOHU31pvBrlVnEmDMyH/ReNna
lUM6ioYXFE9ZFanoMb88CoGYB2SYZx6mLMwaqEu6nvHKxALwR4J7ehJBvgn56OGU/GWAvUZ6KThD
p2zccM/zgSTAELlfblNLvFUKpHNxwo9KpRGmr2d05VF7maq1ObBzgC3BYGhsXY9AhRaqrzeffkwc
vLuFI6J5YcyO5RtJRwuuA7XoaRtbbrBvNxJ5E1tslUpgmTQigcsAA8MIw3ttqvigH20ZX9+lRhv7
wxgRRBV+zP30OtMDgI2Ec7VOirqo4gNVlbQEhgTDKnSLRMQ6wX8s3qJcI93o2v7d7ZcnauqNKp9g
7GSqfnRoFhmV1OzP4LvKbt/js7GApMV7Jem3dcKkUWpZbCGfFmSFdqdqmqg/Of/e0i/EhTxrrfub
+wixTs+A1/7VoLUz/4qD1Rq5b2B/OdOPvBQnRUZXXIMg6qIRkNcBPWQ9nWbdcUExTbJIZb0ZSNZY
FGlh1f0A/Usm+xFrtdTJr4L3YjY2qfJsh5dNIquLZZGusyCD1PELGLm8ZCGM4HqY1y4vRMn5MAkI
ArBLs0VKEM0tRSklxTomHz1jNqTq1rpIdqvmISaAYAUUre6zkMbQq/LfqQyWEbMPAWfjTvvKOKpm
rluOJUiMWqYmM+y4MogCBCWnr4Q5dja1K4wVQHB2G2JXl1SPbhVBycR0Qxp2GfKZYAvgc5uobCIo
MfuVa+mwpOuxa6bF9Gl8xW5Jb+vD9bUvzbW8/m8yxGvVdymlFK0m7VvKZwobWV9nO8KaUBVoJdSl
LV2mz83vhJ/naQJNnNLnH0AC/PtdM/kx3xOb/7LaktNsc/5BFv0/XrCCw+DDb6bGhPa8IwzmnjaH
Tbq2OM457m948RbsFMYF3cOBzBIGqxbA++5HCCzkNGE9PgwTD4uemWfgkAi20oHxNbzEGYpzgOW1
hXzUP79bzm6F/yUkunsnySlUSrCfndkMrys2lswsFuvtEe50GSq8SO6eKekaB89IfqMB4D5cKT07
iYN2RDMGzTijRCjZfeHDhkMXQPmR9zhOxqX+J/1gUos3dYKo2kicLIiQ+O74O7JW5RUXq2MCY5QX
EoTLQIE6CTY4hH3BH+tzVfWH3uvzn6T9uCdE5jnSQtyA0KxRjdqTIqe2r8jX0lzzUN0yUivayUUJ
WOZt/G/UfSeVK0C5sF9Q7ruZFLh8yR/r+ecf1crIT5Nejr6gWvRy2xDRi4PEgjg5OMOUkmSxe6sJ
D5a/3/iXieqbP6ts3i20u7BCHJjk30u1RyTPzGeBh33XP2BEdypw02zu6/xZSw/SkpBUFtzpYgcm
ru6Nb+yuIEDjlyfPJZ8aCwlXrWaMjrcx3f824oY6nZtYLwVT0T5vS9FDvWefuBE3v/Hd+5zlE8u4
ZNR5cQI4z8UwbH1jP5VxhxbX/SmygPZdQ6G1H0tTQKEg0KZzKkdyEDQieezLxKtBk+Pa59YXN1Gc
VsNFpCIeQbfHuEEPi3MgD75QNqUP04DBwtcsPss/FwE6WZiQXWtKTo9dWZgCRYSSnHkEMH572Vas
kWSND8E06MVECqmyATjmWoityyMBvhdF1m5VCeG49Nea6WbX/HFKxMgQsZaDujSeNiqbUGnLArlM
dMS2z+cH1lQ+F+hTd8q7ON/T9PowBuMkUJ0Lu+8ogQwdkZOkRYAGX6ZsZFN0GYfrKDrDwrdejbPL
VksElTyjehx+kwKhreTmM0FFpw3uAvkwTEBsjKZkBiAnxFsURcVd/QgXNpcTlPAc2XXw56Lts+Ht
ERwYDo2435toDwkICQzpyfGcWKDKubENYURMQ5KQp32M0m0avAB200lnAEg6swPG0t5xi8PT5cON
isAO5y+94cPSa9MoeSlkuABsV3m0VgkDi5Z36w2tASxh69DFTBDbAu0t8ifWIzwjBDz0CELgdylq
MZMvpuoeFXGppfnR9rdgTvunMzGucF+pIgzYWV+cU39G5Jx6vA0zjdWjLd+ULLoSp7VDeKP8vcZH
Zm/UiW20K1hXxv0dNSMh0cPQtezIfzu75DIQq8mzfZNRADYX4aBfb13v7HOrMwwtGEmrdVpMuLgs
7bXPN1pZqotfBqnpW4GRXa9vrWCHdIQy90g0BpllrKtiNid7zi5+OqGX1rA0o/K6jqOMGuvXipH8
lvLzqlgRQ7YlDminsCNnNGy5/8AEWTnSo9vWDZYubl8QCVCqfHGjrEw7803wzLIWejXIlPujKm9v
Xnxc1YvFlkU7azda16t49lVVzcjgb+XB9sgJRyS7bg3Jq8mZMiF4CYEzizW6ioyJU11xEr/8F515
rbRmDOZwqGkTDIBZXSGcyJEQ66FJf9FGnv+9LXKtLV/j6U44IOimRdduEMdOVpBQuAaCDjwtg5Bd
kehvf82WymLLdBJPOo2LEdx1ZLARwschTazJxbG94HiqTEMkVwjfcbWjViuxrERJ3WxjXegKO5it
2rFPq7WXjKE5Oor3mXR3cJQpGY38qpeOJhU70jbD87QtVqK9Gh7UUYYiBQk4vdyXZmTAC55N5a/v
uR51rtqkaet1obiBexzgSohMtl5BcVbtAi/FBdy16d11P3HKz/Jy/Dur57Tk9/ejZ1Jr+pJXhUXJ
+25q1+4FknqynADLoJCCb8QBUWLCGTDaWapZB02Wro4HEiQFxorzskBSm6ItD7J9Z/CsSejhCfhg
eXTpPr+S9517FR3PIncNcHVVmSg293/oEsPrN2sBPNDideQ9dIjbkb+/GmaveL8S4N1rTbetbXU9
Zgc3uMyFQVXIrnIHHQicF8qZUs5tP3WBullHl5SZpMgY5mjY5PXODNWTsDfEmubsMze+/855tjJj
agaedag1mv0LW+fqoZbH5GGGPtppo4Vlc5kvhptQ4N0k9KRrqdaAUPJc3cHDvWvFumN2cxG8CjXr
cDl1ZKyodd5PrRdurjKSuMj1et3GCS5/8rmdzZpdL0PY9pmrvbNTTltzADl7WMS22DJqn/r0+sM+
hYd6fe+K/2xl7ZqEvtyZ2DoCvc+KcqfCyezi+NmjMFQ70DAr5ZLW+M677yynZ7G+xvxLd/svpLpL
vtRQKUg6iZIpOujfNYMBV+k3Scz3bInMvBlYa8BiEoVI1/sqbq5FhzWdlRgo16TTboaTxoZUFp8w
YlBv+Dna1eN9vemh7DsZVD2i9saRhqNqbfTTRC8xGbtpOnDZ+IN/6E0VdwsTLCFsxy64tk9tBd0a
gPLwRzPDiNdCMO6GOfgtH5QLTaXDpr5t43zo0Fg5VndIQW/is53WTOkreYQNsnidn5rhst28w4OS
E8BXrJa4jKVQyync+NCaFLpgX5PkY/ZlaHMmBXUJgg/aOOT6eZUCVR5KCF/covw+yRvLG1mlfFtq
nxf/owQP8dSdaT9XxiFcdPBtOT8qTVG2ltYJJwVAQKflMlW+8X+OuFmCTJpnSHt/B8a50pjTCSKr
51ROmQuHm11CGBcFYKqR80BB02t7Fw7vwWKV7JwhjuDUpLYPsmRxvlnpoViKA6fmt21pdq/jKequ
ebSooBJKBhuPtwvbv+T8RlWhsA2BsQXKuFaXi/NYZMK+F5OhMMlaBfFapXZEcfMOrClfd4/R0YrR
nmWrlvLWCxMyxqcfPqljPj4Lw0/ncKXDNMKxa2Z0QAMLuAO9yBEXYlV9bjiuz2zdy3ulso9HkbIg
b0ChyBznvggpouVzA7kqwcT6+YY5lbdaTDjA2aXckdo/k6L7UQYnFeRmIZ9Ezsrqy/nHNgLbK7I5
cBAQ+PEjZFBuE/CBQlqYVWnsZt/ulg8H2Xa9613qFHGCBv1aRNFd1FCzDSS0k6Fsd8slj5CAiKOs
UBUBpRDllvAGX6NKjpmEbgPVhrgRGVzyyKjkqJBCoPtZoTrWZTBj8vweepem8KhjJ6bjl+DvqAXo
xprF2bNxSJRDHqe+EK1tuvD8OeoifA6pe+1TPKQXOPvg7an4tS0GtYZGZuXjTLa2phVudG0JcYLR
6NKS0bOo/se7M1mKdFfgLnRsROJyFyIcSaM4vQ0//c5TNuSuT6NVOZxIO6XkwyvwT4T11QP83QEZ
hLND4YbpR5YeifYbjxupE3nnLZoRCBmpTWGYMiTFmSc7j9ezsmuH1V4bgR4qHMOLA5CXFU/HF+mh
bs18ovsNGK1xDe6c1Aq8REMsV5eGhrUJylOTgZHKVwNodu2wZaooxnmaZu4KQLfWyLa9Vpo3X3vj
xXr24NhTCxQ7+27WG7VWtJsYha4j6izNbWqs0n4lu+HOLT1YT2+gdr+zd0wsmnODMMiEcvj3s3SP
b2nDzDLTzs8c6AUZjx2xkyv4XfrK4q3iUGPjPDv5AKkXKIw57UIzCIfks8Oyrq+SZ658qHSeavek
E4gkZm7UDNCK0l2xwemB/IkBYIEk665oGAT3/YKYtaNf6huXmBCqeSSL8eAl8DiaRJPhcyqChwDY
2aRcr/A3eo6B5AS0zXBkJB4taBUrjwVUJKkfCMEzVLbV+NzrBIEJcAMtbnaIERaiDLK15lki5OKL
S/nLFp3XlrhY+zt/+pGBaKeC/44lOvfMXu7RkPHpZwxdEkEaJFKBormrvhnsWERAcNWXuR/YHrGC
UX/t2GLaYDnq0hTV9fXTrFjEbJUWxMJ+WleACJrje2weZytOXOTSYfnmUmKL3qolzSjqSvtxyaHJ
C4rbDEsCihVElrgu0XCJJLHfBwuvQTUfNJZF6Lf6DlZ05x1SL0PbNLKV+IEK+vqneYjWZtqpReTw
x1/C/heRRMVwSoFi2L1CYCi5DdLqwiefYDdbrqojlDok4cUO2He4yF6dZvXUi3jc68c0NigkQiZ2
rJB46ZYRtc8mr7i4APkxWJErwyXejbGeo8R/PbkDuLv5QMc5zQIpkSwSLmzgZDvWpGmo/bUdQbkp
zuolXqVEF12SPAUiIeuZSD4gzWoDbsECf1gcV1Zftj3VpU1k6DBa2t7BDE8GCxX2LxZw5AthX6Hl
uwv9AoYBC5nvjwKDuhG2dwHJCC7snLlNxwdPCdzLeCJhCyvq0G3O6U+ly564tG56q9L6+DAqWsvO
rdEcwCwzeDUrVrZ5IGeL7zAgALqC4F68X3AeyJKqUyc2NjK1ONzpfRJEyTKafIF9Z9MPPJDQU0+p
eHMpnqmksVizRRAIKRdOl9ne4zfueaSvrW36CUtJ1LNsQEISbFNpHgE3+XGDb2GwUtkQJM2IEmE/
Jc0FYyolBDuwdnwja9epBVfhmyeYapTy7lKZUJrqgt0e/XgezOSJ7GhtuG86czhmOPnLBf3nAuxt
LODExH66l1xk9L4iQblppgeQZ9luVPXFIBCKxXjoBkVHx3bR7z+8UNIQoOfsdFN/IUnyrVwrl+q+
CnTPg7jeBkLHq7TNg8oMY9fvgYGDZL7yv1WDLN/QLbG2ndMz22EOUDiSE9dEYta8Z1jBpb6g5hmf
9NlXRl/wOJBXO0SFMvJMrpZPGutoAyDnblALJ6n6nrwhVElxh4o/Sb5FJKopMoeCBeopWxqA/ljq
X5WkvEieh7CxZRKXWXTeBI7wQDnpHrd6DZiUzPaClrfULP57Pkjm1GpWY+rsS8Fbm8sOXdNmhaLZ
4ekQA5YxOmPNBGDJA52EC0htaWaVFngEIFBCtgoq0c70BRzhKp8mwYIa53BgLxJoXUrO6qYtRYzQ
E3H+n5yZgzFiw7HlrDb+aio99kO6efoZ3ToAcUGWJ7m3Ss1R29r8NbctWEPJRgdfXoSUYJX9DNb9
Ey1NzDCVxFtJdkVqUu4VjE2hpHeXXzQso38pEXSk68rQY1T9+eIkpVh5y0YSuoQxLAa2ePXBL6Tl
3nOq9wrQKWN1X/O1nrANoWrnjBb3XEIDmj68TazM6n2Isa02DP/GHPr9PCeNw/8KZdJ1iO07CPMz
5dqr9f47cnmYH1Yk9eQdnRYDvp+7UmtFNKc+SDI26M4WBYwgvuKHK6xiBJzQlnXQ+6YopSZGtaFZ
Wuu9xY8c1ggKMFY0aRq4wftXCySbA9qOVArbbiYSCVAZ89pnVeuksWUJ86GC4FfrMv0j1qUOjuXK
rqb/LtzlbgapimAOvol+4Ona4uEDrgfoGmEF21O+tMrj08pk81wCsgb/1r1ZLkmCOW3ikZONLPn8
JhmnXrJ0r+jwNgipVghxqvVCznh8YnyS24C6QgFi11Rcu6J523gA8a7BlA6Rw3EmiL68H+k6UkYa
D9RAqtzbYkswCmLWGj13L/gMHa9alphaSsxyOmzqtK1dqVi9aPbgGBmITebcSBwomnnIpVuc7A+i
ZvfSlDATtUgN52yb3aEzdR1slHk0WeHNaC2arSIF3lUl4dz2yWZgIR1n6Yw9UyvBL18AB3zn++EB
oyQ3dYJFGBC0Zw0bl/JHM7haV+NmQp/vFgn+ZUuMHV0xktkjUR5AFFVoMWXhEnqGM/AfhX7SxO00
naI1WCRGWy5I5/I790x7/ZSw1xSVAOg+Z4V6MzjaFk91slGsG0hP6A1Jrj36hok1dttjC54pDaDY
VPBiM0nmjxIyRPQ7V6FdS2MPFkE4C5uctplnvI1YOMB4uBuUvyz8CZQysG6SYm/9UssiciW41pcR
/DQtXhuhVIIi1L1t45cgDVv/ce3QnX1JaK5PN6teU7sbiPNZMXdCbxH2wPChkIwgd0fr4xi9Ynli
XQ7AWE4Ed2NX1nVbFjM8hErOM/j/fJqtZl7uth+Oi4jgpe2qQQt8NgxYKo3xlA5s/Ku8XjgPO4Im
H5SYYgOvIHXC3B3Ph79o2pcrV6TLnCOOruoV/93u4l5pXgxNNYqadHCoflrVFkqfHmyg0kgPnQAT
VmxTqtB4PnDuVVzvXY1q3hcB50Gi4W2LDcjcJ9Z6HsEKgl/5sv/Mvq+lXSg+824o/emyFGqvUPda
hRezlJbkPa9iu2Ko82XNlKfCMKLPPYYFUeLJRHmmcKHQ4tZ2saBscEJ/slN4iKVfkZuJb+SHA8YJ
ZE06H8Fq0CT4mG6mrXuoAJ4mcc06A8vOwaKSCfk7/yJi8SHrKiH8/a5eHH/MmhqVBdu+s9nUCjwW
D0j6HfY7dA+9tZK9WL5Cn/1yVRGNmw4w+YMMWkaiA8OymSpbrwnX6hWoLSwIxTyBVj2S0btVko0/
9mTUhfVw5L6vHnotTD7sMt60KgRNVxnobRZY3JGZYWIMCft4S9VBVNDB9cCn4dTh/kdRf7t7Au//
0JYlqXldY/1a/CckyShHg6xkKLW3oYa0A+CfqZn9badh9qvMF8OTEgVAMDQA/e3YWT1kYPtiumyR
Hh1NryQhfuWdQRhZfLJrDWaeNrll+QossmNjyCRkxn68dXKgsde9MA9YGiSr23OFA4N84/E3V93x
s6WIIv4m7rTkzCNN4xuCNFGkjdthU5W2vNysfASBgip7dA9h24SGGBMiH87v3wCovR/n7u+j0slm
qMFdUyjS6I6iMc+KQcIUxpS32TKIJJzfF2Vdw/XRNjmDMWb54wgcPuICH35+I/p5LapTZbTE41HW
ih7Fp0ei941KkH5zVtj4sllgHpBwRLZSJaAnAUMZhhOS4wq+VoqA40lWkps4CJV5mRO1VXRQNXkp
G+Uk4xy2M7H7IQ9ZzuaOPodcwBxjCNX90+JkNgpLkDBBAaoETAKtMWP0RrLyOXi263M6tPyAK+/x
PAewnjOuiZpbBRJdGr6d9398QRPxSmaylX/Rd/BaIiQSgIEX1wNiYqV0cVMsQs6vIL7PZOgp1Lqj
Zh+s5vaVKSRGl+P6V9ClgiYabbePtlXXjAGWq+0IQ64pMgFbcvQVaD7X2QT19j6WW5YXWjag05tC
kF7GqtXzMl+qotxm/sV4ETfGBKdGlarjwHXmJu8sqCVTfMIUGRKxuL/V0qw6425FlgGwei4W+or0
i1zfNA6QcDc2GkW8jLMhgQAJcjnBIgmb31GpkSzsz206HYtPEXe1hF8XkpkuCVxY3bdHtaYcgrG7
M+W2VCBUV3ESRY2zVXheylXgA6cU9wSatfBBj0vmvDfytqYZNMa/XqGzj3iS9bUUYfVESZLcpwNz
R8XveCNCB6paMl1T4ssHE/+ZbzDp16GN4YM4jSmTrESk2t6n+vXL8aSNtQ+7JberJTKUQ5USjnAC
SRgakAoU8cYM3eRc3il/CT95FtkqG3TIsX6nKVHhdEgFkAt9OZnR9VlTUQ1L4UaGQchIhmqYv0aS
/Ctp/b2KRCMKDOyLNCtWJHtN/oc6dSVJhqJY61rUVrQkOuiF1KBHztq27HQ5JukUepy9wm0zTTNA
CmGhF0pbKSHgRU854xUnYsVpG+XUv5+18zGecRlC7lDHf9R7A4ufr2pr5bqT6EDXTe24FBrtqedd
3/wTc7gkV3N2VwfvXxcIH1HZc+h5BM/0Ow2+Pr/sEXZe5Y0Gg+tsUsej1kqLy/2Wx5o/+duEticu
FAbrNvpvHe9YUXdSFvo1j52QCDn73MNbts8XlB+xfP3063E/uyKiXn49Twtf+e2OLDhD/C3uvI03
1Jx8iAr4c9CSQqdcD/ufTihPQYbgeJ2qrL00OZDudPMsqks6WR3zrSYT5lUwbTdj+wZDsQauK7W1
mOKNvaKSvGHIapmhckZxbB/PHRtELSUic4Onf3Rfnc2MtQKRF58ZZeexgHDA5SYZBnK/tL4EVSwb
7yyt1S10RnNoqubCHGgJPpwOdjZkjrVnbSxtY/jeWJ7rWufA8+gJE8Xkd4b31gqHlqYwPFVjUoIV
KUkOsAJewkph2DjTq0sB7ygrC4LlUezvn2qfMkmPVwj5BgTzuPKx4Ln8ITKNbXAkTXGeEd994CvX
6ug/DhAnBkEwy2RsnJ+OyQ1J9u413sqbDLUUDw2TvfyAdmJwuvYqdR5OYuy/6Cwjk5HlN1nRK9k4
MramrFP26awHRRbwhhTgkcTh7OGvF26AXc2AoVg7b7DL/Cbr9MCQVhKYYOVk/kRxlY55ntCJA2+Y
a3YXVC3qaawwnCnFYwH+2oLJXMzNXpv+nNZiFnbT5Py6qIaK6lLP4bwTZ20lYSNj3HJ9NEUE52NG
gSQIBhBvLM94ndncg957g3VT11/M/pFcaUTVQJWNz7QnLX0RTc/WUO2a2FNKmrpRn6Z03xO4F9g1
OfXRjIoJvy11ZIf7rn41O/6jnb50WfmdG8aDFIvd73yAdDyw+hGShBQLdna+CvzKsNdQNBComyyJ
uxhiQdMnVbbFuyc6B9DsXkM5Iu/WyR/IRXHzIvTgFdO1A9DaQwluCfZE5N4GSOENv6enLMNFUjJ9
1jfHUBnlZifA3sWfLFVFkHjz08zjMRcT2kXjZUXDImZ8jdz594GY75kYRasCNM5i8vN7N7uFkxPj
zuxSp/9mqmEGCv2kqQ+SFzgHc70gmntOIQ0GcZU0ixDELmoZ5iWZL9X0mKCSLI3rS7rpIknnQvCs
TQSY6zx+za7eWEGSJ7CkOCmGQc6wZf6YLWBu5Z5kVtg2i9W0dO6hgXOjhytTtkKXSXuc3nd8Vrqg
ZF6AX0GkP71GI86KLLiZP8O7L2K02fmcEyM2dx7GN7hv4WEJMB1auzkAOBLaB6aXsWYXf5aontmM
SJk4tXhsMXdSnQGlFTyPD3glm6c3/QQyrosYdd46Xf29+TmGy8m/1NppBLso94/nK8yjUULYSuTy
N4rE7cqAlzX2p6F6l/qNsZli/svYpiw0qXfKbAAFem4VbEQ9ER+r2cFywtRXTD+aQ5UYPsPAJlaD
ga01RmAHI2Sjr8M/aaH5baGvCO3LrU+17L1Ve0GxZkPqsmPazBCih1PCSNoyxgQ3dPwoMO8c8Uqu
dE12fKOC77Y5eHOjoppTUsM5jc1t9j/F4jnogI+hEucQ6xsU5Os0aDI6rJMT9RHytoOAkkroaG0o
Yhf6DLhq7bmmXKIj3j83TGw2k6MfmwlIqIZlVVUk9UpVPj87M8B+gKY1+luvPGfmFIPaDabVlzl/
xYWeilb8IiT+BpSaQZEOcSiG3bQU64DYhTYbzCFlICwPjUmXc+T2+0u3DQXf6PMjtuM93Qd1es4I
WTtKdWosr+dtCCPjPpLwD48P9XWHXwiVWP3iriIM9BpFxRW1+ozPcezhcOERUvatr4Foe5l0OG3b
aBuc7YCZm+28MCjDkEbnDcEIeqJ5GMNdD3wT9B9vv/zHr7mwZtJ7EAN5oGTDYXaqdVMzd3e9PJXX
WERfUBj0thxevOv9KHbyGHvBnC/SrX6DPph88A+kJOrropiIYD7HdEKEARE2V/E37Wu9dOP/bg8s
Ggk2AfM1bEafh6FBr/5gz3AhiFIlORijImB1ha6lr0ahSWvBSAm2G8NVO6z1i8Jnr0qcKdZ4kamK
ou28TpN1zV/iDv6UYk7qPHT3AMFynryky+JVewFoWvGRYHM692c/24yrG/naKMkwEPJeVdUT5UWq
PT1Yh1r0zTXicLFqAPEA97fc3t4pMpDQaZAtPZoBBWBmAL0gcuI+uue8Z6xCD2loiqbV0JxyhZAy
fKo9zjbYgHyUmmn/BMZs8IMBLnzsX6EeRXbmEfEVHmbwwZ8i/jEadDKyiBOfckiBpUmcm0Jm72kp
GyJ/dW74GKtfcjVprMn54cyx+tzp3xtGonIoLYXtNcABDILmz7Hsppj1lCf+2fVgc37CznNAy79a
kh1nckY3cEU/iJop8nZyot2WYAL8SsS2Va7fqpuP0I5shdEarm4TTfyhE564Rz3cMZCd9WMrxPLY
euFCxY+JTUbHyZeMfHhsBOwLC1Bsfhtx0K9EF5WH9LufwbOHN2unraW+YzNWGGJVw3UEvk9iVLIq
ABb9N+2PtfXPHS/5iweOmttBORCZ/T/vdSS6zsmRz5j9sbn3Ej3Kf7tezhP178l84bwqHhThfcGP
Jbb9dm2xOGVo3n8CwTf3kwGKOJEWTVTnjrhl64P1gFICR51Y0MAaM6HCjCTRCKc++I5XWv4g9Nm2
aqQHBdS6IY45MbHbqUHvQrwrLt1/CY7VbFXku3otFNJCh4USjOznhmD+zKYyfn+XBjTimxGh0dxj
IrFcIMt3EUzSiXViY55r2bS7zrlBua48QNUZhr/M17hQ7KV9FroUNxBqlXbGHIMkqerXK0A7aABf
k5EhHr41O3qSnQHgzwOd7FdsM2KgouCSidvHWIYYcfrPLMOlbJEaKYvWTaDhzcjow+AQ4p7KbB6q
e+sfl+a8mAeKuVBS/MmfLQEjNZ7FhAt7/RqnzOUtFdiUcHNrfMai3Khkzi37ECMTu0QIqZvPG6WY
z9KnNBXsjceRp6wvnAJ7Rr78KmfBy2MBVmFv/N6yO+Izb08rjWo4V71dMl5YEKTuiSrbU0sAlEo6
Wzgxir0c05AFo+J/bIlCP4LWnV5MMCLQ4qdkBe6j/mqFtOWAsNIzAfK2Ddq9812jHXctbgGgZxPI
L8tKKsNH/itqS0McH5QQLunEjmoe2FzObPc0LK71HBSyHjVWfUmFhSCQiZD0ndVwQ13qEAkGyyFa
y6GOLhG+flFXNlQwIUGWfBDrsBeg1bqKUBWeV8KiJH5bD3UvGoRXy9Shpps79XLH8k3LISFw8yoQ
9m8BNkW339xsHA8FZtePnJJzjWzL6o8CsOUNqJh6+BCZm/Cci0Cw7XZcxM1JXUaR86mJSzfqavoC
200LHNzA/n3nBRekY5ZGbIrIyynZjdrUF1f1SO/+WjpAaGIJEk7/HpAi6LssjAbXduYSFCgh4/+c
4MFkRXY5KOiXp6Q3+Ly/HK33L6XU5ajrS8DDXmkmqH3O7vq9QAVwML1xOhTLBgrrv9DPrh2kgnVX
qAAVim3wwhbKqdb1mZBkIHK+3uGKDKjEYNTLRmThwhMi7x2Cysi1YwmHD3tA30+AN0FZwDMOMW3F
Sp33f/W6FBDzmOgQYoRedww4nsTVcsoIjxO8va85InpEQVis9J7cG6cdytpBuwEdt698lcJcSstO
K29HSp6qNxUDugaBbWWkWwG4dZXbsvyFtPG/JFkd0ewlHQwAGfltSqN6wkmxIwXenDMyy1kG2K2Y
fuiBJepo/9OYb3gtceUPjV46b+v9JvWbJ7de9+HcmwruLvsHPdGAcAFJxuiI7jj28WBvL13xuvLH
VGKCU9BB00ZienmU7kOgulB8oBwsaHJVLVuzJJruDj1XNZvlmQaOMzg2UAM/LehHEkAxKaIXP0kV
1QUeCrWWTYy2BKRthnnpiHF4V2uWbBPuWQRtnl+fbyToWCIRzjxoy5G158W1dnOASxFKVmhKjWH0
/C76HVglGlIiqfebt+Hdr+eXmCbziOdMofHS7w1vSCNsKr6G4D3J/FU2co69ixG8jo5Bm56Bx57b
MgU30o1Ap4RfQp7ON5EzE56qFQPhurl3+sycaFLRDaGuUnLcgidkRlLFhYCP/SsQfM8cCqeQZzSi
QON9VQREbMkrtWyPzaHVQpX4N0Uww2mauovcam9B3v+J7WamPE2c1WIRgiJMlvAemGuTQIwZZsGs
ftqYuq2AiLiw+3GElvKWDndrjctnmFWJCELARQUqiCMR7TxssVwoqhFz7XgFO7YHxBAP1TmOpxkv
u03NGoUPTUTY6kIQoajgYZ478cKg98ivZPK8keT647ShrlAursE9UGrMD1RFs4QTLutosgAA/x57
MFfiqbUFzNccFg65RypbcT+Im/fNx5/E2F4SWIbwFV4phkGctcKx7X2H36DvMtqZHh/vhoz195QV
MsaiCi9Kt/UqCNeWHTUsT7fu9PTiIhe38uHZnyWV8VmbrFL8WzSwdmnKB8qBzSk+Ii+Xno42iH1b
mMWsStDkKN4q9BRaumOsX01LCsWuQH/2PlWBg6d03pV668V8DTKtW7mb7VbUg5H1cGvfF+0sAtyX
VPFETvV9o13I+rxV2O5FXlP9jZC0gWlLMKq0bNPcAZN9ygnVVSjbLFisecRV/aoonfHkUdB51wRi
wW4+Hh7TZfAkLdqOzD3eyaCJmYznt32a7DBwtPaieldvCxoJb7qBGFxwY9ef06V2cnCqqUE0uSqk
NZ96q8yzM/Em0B1yNJZZ9eJhzgnf6EJhKrB4yjC4uyMH+FCX3F0Nd+2YrwghROSkrg2v/KBca34V
0FkiWYJJOXliaPFwz9M80rm7DtdHPtW86q6B8LQMCKrNau1qjJPTECSsLKUh/W3tmXBqJO+G/k+b
rOlfLmOYEwNW/si1fY/vZ0ib8p76hIt3U0N4WPastG8MqjDOyQTvZiQWhp/nqb1rrhFF8m6BXZKL
NyKlb3eoD1cMfKag8qYqvTGlSs5uFgUAJRj3v7bRtu491xM1Xvd6X9ze/PQGxxNlT+pLQJoXrZ10
W5aH5xBaD2m5pSjwnaKG+cW3JkwPTJ66LuN+cLnKsdZzMOpzefLbBc3wafaUDu2cqq/HWPcCoHhO
4XpeH4po0hi2WC5stiG4AVw9n0grn3wZ808KMqASetYQUnNPNYeSurQR2khHhJhWonMcS9AbWAl0
IJZ2/YecuNNMohPQcxbD4G0S6wXLBYixCjwo2S6lLEUQGkNfxHNi+FV8/VCLrf/qgqdXQJVGuvZy
7tLqgFUgY2Tpa9Ur+XPplSWVo56rSr5AWd0zlzL+Smgl+lXyLsNVXZX8XBdOA0yzX7ntF8TBBoid
UGVlXefbN0hW0B2F2mhXfkIeuwJbFoqMR7vrKOQW5aXqbCzIamMTEb0OLJw1qLPTiW7dt/w0SdBj
tQqSUicNs/ZRbE10TuLXUeXjARJ0r/n1di0N/17L9ZnX/Btg4czL7R5omjJFkRUocEw7MFdBYqMd
M13/z4O5U9uw5TxyCLVvfn+IvrqYmVDYYgfDlOgIAZXHigCBsGX4ElaqvzvrouET9MmzmGVo2QBq
9t0ln889f+DVb7H+vynD+wbDB8kFpTSlyO18/AhsyStU7q1XsHoSAda6l6ESinokIA7n4pasdvPG
wmN+W6M0KgsYtVv33qjy0YRTay6S6zDBiGtFBCtI5GmBBfsdqFb5NgY9hpAg3eUisHLgLwnkavGo
5ICnBqJyDKCh7lbiDr6jd+9oGRqxY5nMnC/YcX7PuikejMrM8uERZ9V2s0KqS4dkrBaoFDp6lF2U
cwSTxHeyxWONxMVRN1gbjQ9J4iQrYCQPWjAY2rTnbIIXMAQ6Bvtm8+8BP1LwwqPPQwGU+0kJCEYH
PWJSUpdE2sGPzwxUGugL1ft2K9jcmAeKcXYkuNJ3GsqmstwMf7N38+LuYHzxL+MeFzKLvBcIBOl/
P7JzShzr7LxE2Jr+34VOqYxOFAhUiebL2alxj6d8zCEvbJwVHEv8QV/+tUvbSMz/QL1kKVNn9vRj
AmJ+RfMjP3CJByOoWm7usUiCpWweIzWnO2wcSduO4O7XqgNCw8Bbw+8f5uzmrWv6ozDAxYHbkIMe
Czf91tbXervfig+vOygoOWVDWD2qb88t5naa9bRJVqRg7AKd1VVY/VtMkODkCkqzhnfdTpzcn/Um
qnlhhkJgJFzChdyedM/3y4l4BO5k3pK+wlqTx8lQ6QU/miL8iVmqBTHRl8uBDpj9QJcndrYKaUxO
7q7D9yWBpOFqmb/uyzypWUPTjnQVl7XSqJozEyIlZ2Sa+xZBrynxiHs1NodZz6tZoqdmL2F4MynM
pWjmy+Kr0cbepqME1rEacfyt25K+znQkl8nzVDhRCeRLsV6VojJWmcscgtPrGTdhSNgPZ/nXr6Be
OZWQ2Eezps3a2N0Nwq1D7YLtblbCYIJNtk0HJTbWspsRnS8fAn1SByiSk2X6RGe33x7a1kvVVX+W
b6zeepVVIuW1gNGjjHyk3xkf/XE0bjGmTL/Nvteb4dE+K8Mj/g6wXxsMWC6QRQpogzWDtAq+kdg4
b/2YFDTnlTdKfh9Me73Jgph6EaBroY0hZw/FBe7E+tro0/qY63eM7XaDv3JqYwinca8NNcuwzNpw
9suswtcBCH96DMKNscRenuLdFG5vI1IoBNR7dQXsrEho5PscfAP3J7L+Ltz9bYf0s6EpAVM9hM4A
+5wIvq3vOuwDinDqNtoH8rNo2D2MiHOdFqEe1/ab/aOyyMVQD3BABmHYG6OeZdRgZbQVC+zkqn6E
03IQ0spPXWitMUBR3yA0OomAgsZyWMO/wo2sL77TUNZRCm/2cKHtF9y843BUDBKrPFS7rZuln1kz
SIrhi3NkT4qbAFlrmCQd2zOaIRW81rwlEY8YWTdr/E+2lZMHJVTxOOFtAwU5wPmeCWjhY3b+ddHl
lc9uWyPiQ2ocGdUJIbZjgHozrFHCcsecTGGNUUYhsnpdXcHXzSdee/bVn027s9PQV3sNLs8T4iUM
lHPF1VgnYaNjXbLed1a/Q6/dICKC7h4TmdU/2B0NMFVfb3benmeS6DN5KvedmOLdkEFmivf3G3dC
L1ySB8Dhax5fB75msG1D+Osc5wNo5rPuuFnaqlxbSN3+EDkjgw75XiZdVn2ZanthZZKf6SIQZlfn
DhVLoSMQN6bXeE7A7Ycjr7+QO1Qypad3UG2uiQIAInl5bcxXcJpVJmv5NKCkQMLaaA7hPuBBm2u8
TYLOzNdvx9yn2UJ/MiQzEn+BfqHeVKaxMMrt+lAqRcDeATZyW0JuL35JU20ySIHvUjNUlmvNoyZi
FVJlGp3PS4XmjMq3JooXuU6UGJKSmN9ryEzyvcu8M3Xw8o5XP24Ps5k+a1eUc9hWG2ivyBySwIXd
W0cYqvE1VFohVb7hGTpkn8cpuFJ3T9jM/CZnEHIpIS40at0INlcWC0QN9tNobMNKoI/vIKIF/bEf
PUWeh5l6TWao0AWxlxzTL7vPeXv1HGMpGlgIvTh0VbZhFTXh9Az8HqITRk+H+sALnVys21XLk1nw
AINMisk7q/52Cqwgwo0+0vJ55Myl1x4m9rCbTtpftADrKVZKJFvUQ1vve1pTA0nJ33lLv6AG8pyv
GlWwn6zGbqoEGOcbZDG6jFu+7807cxJB3/bXoQpupwTYAemfGfjBzIm5m3oR5unIkp0bmvd4DbgH
XMprQx4lzZIXUbCM2k5jvCQNQ5i25RfZVGWlOL+8zMMBSlUAofj7RPjBPmJepaSKoOLoxaY5j4Ak
FXysbSwwOR605JrpN4fjM9i6rOD+BZXYV51fUtY4aomC2viN/5SigpAJKJlcGl4U0kMmB6ha/jZj
T4ZjHcW1ugmITByC11gOy9OruAzsuwI9AOUGHqAuq7K21eWQlLo9aU3zRe84nA2fsE8At2Hr+vGe
12cExduGy3YLh26jgzqNclH8QpNhymZJRa/PGWNVj0zGfpazS8nV5GvITuhDfxqDnxJKGy9dI3S+
Qd3dcmrU+lUzh2jd5qt1tNr5NxQzufNxojKbMrXN4t8FuIfKIQCyO/EPppTLhIEwnGLSDVCg6bJz
jfLj+/8Qtrdu6C0u/6wNCpjPag2JYn0uGaUOFYR11/R7hfO2dSZCU+YZjX5iAVzd2jO1iNgUhKJF
nlMjdNSptDXgDMPJKgiZHZCCRu4QxkiUxQYHPGYS0lk/9Omx2/6aBO5OCB1kl7zTwmy1o1ir3qAM
O+LR17qdDHxT5A0K2hqq23jdnE1iGJSLFHJ3oHc4mjiUvfggFIkCPpVIe162PszNOg+1QePfikfE
vwjPxDA4j3H5wr0kUxlgz9PqJR1RyYq02BUsW6nOOuwcA0g/jXVUEebwR45euE5MSz3+SfJhY+R/
qbb0Z8imMjPITdbHXzyLL5ME7iyEgfp/NSAC+JLRclLdV6El8r4K0UY1n+RAb8OI6TqskU7LmXKr
Zw25wkrixyzwkHf0HsljxMVvYwkdhpowrxBqiXMFilC8feaXOYcQ+BKAxjoXpyncxzERyX2AZV9P
jgVW7tbykck8z4Kn7DpW/udZWRHds/I/K1HEXCPxYWLlW80K16l6vl7+QwrDWdXHFECxhORrVQAS
9GFKtS4z1B4msDXBVdEoGdUAcMei1p4pYcj7dgraiSMDpZnfFGxfGdZYIHOPXn9vSoYxcl7/qMEe
bqz/SK+16lubc5Jb5FMWZzZbxK0ZwfEp++ub4UFkSFRjNtkktkc/SaarOH6wLNFk7VE1cYUcM5CB
IqR8Cos37ypcpwyxS35vocqsGkHls3Fxgf1f0tZiP8axlijecVO+6ggrvd7vKbL6OZ2yd5zSy+9a
OWXsAooM7SfKT2dnS41o/mSLi5pR517TUmis68qVbNGRLOVhw7qQIia2hcxH5ePkwr7ffgdnOnVS
w5oU0K8ZVOVR6UZViatH8JpZtWoqrCsGzZ58HB197SGsyFg6lMV/laC282Sp9gpxCrRq+znhorjP
Lbphotaer/aJzeTTEjp9cad4PmPh4HHRR7ePCgyi/f9MUVYKr8FL69vr4RdL/W2jH8ZHSEiWGbAM
6gBbyuFU07yGnb9sE3YdlLGMm8lpKRB62xnz9gxj0sskeGAjpdLDFjf5QeuyJ7M7mA86lg+kncli
UmlIdRg5dAd9Uk3x+IryRzF6duzvJwGCztjHxRUd69OWXWODRPCJ8jF4Z86a4fXwIb1ZUWaUG05E
L2Cfoe4XY8vXbU2C801vB+vN/hfdOQ5mvYfgUFgFaaeJh67rm9zbZ0AO5EB9U3inlVMi2mg38lOQ
btbbCeVEAaclWVL7YJnxzYmKuo+wpyyaGn98rMdUbtq4I6hDmUfBSjYb5wzjDrGYLcVf/m1nGFC4
KnFoynWTIMmnvAZpaDKjtJXmKlLLZsBT2aJPmjP75p0hmEogFDBFX8qKg0gYnVKkIMx5TOq7WaBy
AJ7EDsYG1R+twmKukcQrW+cesSh484+FyFW1nVAxGyGIrBHgP0F4fZ1cmb7NTCUQrh46i1up1zuZ
Wd0HFPQMxLSKC3I3RdBhPsPAMAaXPynoUXNef7GpFDeNPpYiTvWrvzFEGn8rSqgn6r04rHN7LDur
3Mp9SKNOK0+X3d/F36INcSe6BG6kLUuDCl33ZTPctwjdC6f5SsedZ2z45yHw80qg54MpxJ93Uj35
T91rj6ClrmgEizcWiXmEpBx4W9zC72UMNS3GUv/Gxub+7rm8vawWChWc/lG1O0ctLdSn5Fjbp18q
ofKpd9sgdL3EtGfCiEmRfgB9bLLSlb/taFJYiW088/c4cItU0yyRlG/rMM6UIUEwV2lRA42MlglU
T4VqXOmuae1na4V6zdJjqXAs5n8iEGo4qnUBoiA9KQjH1jxpCgkLgwxcstbvMuv5CCeJ7riwu6gJ
fvyTjSLOwoq4iRqUtPSoXqpGXhrtHCWcySdycp2RgBjQVPO+UbdtzdBqPUwfHhmwDr8hWY+yb7WZ
3MwpWwWhYhp52vNp+fLrdw53WUGnxZDDfAyzC2fxmW9pvGXK6VuVRilj7fJtbtM3DP/Nlx6riet3
EbxRyvfN+LtiIfWh43SopeyVqllJ8Y21Uh/iyW+SBjB2ZCvxUINqf4RmWHYvLeycIEBLbrRwtfD+
6WNGVsNDNOCR64P8PHIsjZ4kDdtj+zcu11kJv96F64Mbs0cpi2u0JFZb6SkoKAgtF+gBe6jd3cUp
Ao/y/12WPNoBhSH6uQTzqqMLmemzSQyL+1YsRf4q5iQhAr6+2YkUsKv8Zlhpnt/Gzn3A/d1D0RRJ
iVlreHROpunSUu7H9TEMB6CCSWA0XXtxlbJcvJr3AXaQ18m5THqJUkaKQpE1uMzrzQttKUc9aVI9
uGL3hjNzCck4WKWcfj/PKtT5QUsA51z/GZ24RvJXzvbfFWPLH3BL1YNCGr1V3ET0t8rIaXdYfq3A
Ryt2itBviizQ5nvn245bDBPgrzCqQ+41Hr5EWZ7T99tN++kzawqtNu14zaDNCdBvIHLXoykw3szh
DSk7oGE3IOB0fSB83nQ0Mg66beeB3idn9/uxLmmQDm1V0KqDDBIDU0eL5CrELtzZgTi7Mov4QCQo
PC262h4iU/e/9CYkQb5yzxS4oUW9PnVD/LPZ8YOMxGz8Z1qDK8P0HfOBq1AupfKGGCOKeJoREFh9
tLkfmKHadzg5Ha8kbwuzzRtM9xDnvu3q5Fhvhy4IDmaUqYS/oUb4021uvFFWFW7cItreU8K+Q0WP
vKyc3gRWJEgsFLxiWL/xT13EzZ+YEaKFAxnEVU4IZl+QazLFXZibf7wO0TD1PKMuqn8qAnCVCHQO
iLcpU5PyQrtKapPP7Z5B2AOi/njjN8o8C5UDYUCwdZvnFzQWxJlhUadxzBDiETTutDuc91Em3Utg
+w1PlJlTGxVWd0w3WkneVrtJhgVvltoWIN88BjsS56DMMBkWyYJh36AxHHP+WU1ISY/e79S0kd0m
EZypCeqV2hQ1ExhLGeXzJqcZwhI7xeatFlb48d9/JQphzNGII2PcObM/CIfpJ9You+4aWQfEjuef
COQHTxXSYkiY37iZh7V8uuAdmt7fbvEB2AcPppCc25B0CHYOA0bHD6443V0xFuFBSrnoVtXykWHD
e+HnR3NMd/X8e1ug6c1kzYxjePZNXHIKK7KgoBbh11FFdkYBXB802XITRojljVJ/+SPruP0aCeXv
I2bzQFGjrb82eRT3mxE2om5OwIG3l0LDJECTqLWXPza+VLON98GkfhuwegzIXPTKwm4CQS6ps+Wo
O3Wm6IzXUa1lEdq1WCFonGQsflc65YyMSpNZJeU4rkOVL9v9xjv4/aH62uKvHDiZZPthwKwlrnVE
rH0NA4t+Cw3Gs/6iXXMFfwLp3p0viUtx0gPAANErbs1i0+ZZR7a9jKJx/kEAWr7JSRbcMv09b4zH
Kmc0K8pIlZuerOe1tLZD0Ryq7Rc5Tu7kqqyTcJGAl8j69IkY6Uq4A/FgkV74PjHR8k6J0iN+uvOO
7TdXCgbpP7XwD/fVKdcTKlzMcbJxHQXFalUh11T8GjqTCRnfrzN793BAmup5x0HwEuNmRIXImFzy
5ok2gZEP4x7tmZyy9nadkiQckY3TfABxqJ14E+9zL7Oi/xD0Ioeffs2SGWHuqgc4i7TMD47a6tBl
qIXHYgelmm6OWb4w6YgKX6Mau1W2tgLOR3xJVsxWo+Z665GwBh9WmnQ2swVhRwN7nzEWbCntj7fq
1VqH8+MsH1Vi1FaZ1Lm42JguPdusFCrDTR+F6xx6JlP1krQelneNsPdZmpnNV2gY7FuYQod8xXHJ
IagX4sQyc0l7XZPYN8lkySstIhuwWqkUwU3zBQL8PpZPhCSl0IwHfI+dDrcbPhwn0vmIwHc+4SE4
Tdb5Iqe6Yhcob+JmQLYVA5AV8jUw3xH3UDbDsmXKbuFiCPzoEnS3D584mW6suTB/IrxUUBTaI7x6
a4uEvSuBePYYJzI7ub/gR19/kEitMFpDxYhjHdBxa4Lm5Bzlx0P1vKq2ajM8Z/4LIe5Nbqd+K8FA
bJa9pWV1FcHxuVMRVdg1KUJwv8jVVfSxILvmrSOS6d4xOMS7XTqbFnKpm66V7Ybns/oDrAcSZOx/
J69+STq32x6lLFlgfB8gI1fePyYSIBE2EP20VMEbaLriskq+FiMcA1r7ARqawmU43NfqUR24rBzr
QbHLzCpbAa44m42+uFdtRTSA/D3gMnvrO6M/MTwFBhBsicQZ7C4zZTGrIoRf6P5iJnkR4rF7+Fem
SGoGHJZPcSjtOBB5m1yb4r6Rbc5O0Lgnb3BwPdk5WM5kVvSaxKeNWbUUYVz1PSoya0f0a/pyVczY
zH1j9QjeQR7VbceAGAyLtm/ddjnIZidmsqPk0QX4WSfIUcOwhmVLG/RFGBnH4KIJmrsDXM9S5HJa
JcOLDt7yg5UibjZikQq4yqMD+e6Wmp808aisCrfuh5vgOVOt+jgSGx2Ili9kDZ2rVCi/80f3RLTp
JT8S5HxWbW1ucER9cIT4SwWsnR+pTgEVJ1l+Mg7ROlzQgfPfQQMVa3XfhipwUtgimp6UH+G3TxKy
8kTUbHzRG2n7d29Pc9JQfH6IG9oC1JF5AccOUAc2od2uni6yU8C17mmkB1KXn7k8EjQCVhluJ0EM
wSz5JPaJP1Os7aBDAFiVH5TpToOeujVvzzSgFqiQdt9plzN0W4gdGwyiYDfas4O5VRg2AeA0HEOm
wDLr+2Xcw1p4590AwILiyC3jMpJtrOsKo17gBdEILjeWUfs0E8z6nCOssenjksgp36LOgrXX8J6o
AEeAXpX3bRvSOqovuPP1rmPpqvDKklvbTE3OdhsZW5DWmDLSAuL940ucCJnS8aENzUbtAjS/JlKF
WV78xPylnFlUPj3fXnoWunvUiR+h6BtjItPYyVlTx7MQqX9jls94mR6302JMXc0J3HWLrrZgzdyB
0A/VMuidkC7CdrvGwpV6NBYQdK01ocPw643YvGGFxqMN4fFN8BwPA9XCJ+c+JDRNLJQxRI49Mbj6
bVoEzxE2rsp8hguotzh4WP2D3ZwYUZLQyPYzzeqyJNfuaylYsz1xbsNOrDCy+ibYkupvR3VghKfx
PK0+8eC/A7cPQ6H6e3ghg1GpamZlpvjRT9xFmGadWE9x8uO/Q1BclEjwK9mQc2YtNDg8iKUdMsD+
MgG/bpTTveoD5EffOx+5+eKxPGqLNDGz7op0aQoYMuKZ6ir5lTyYoK5p6iAdnL8K1WH+Ci9IskZt
1ujOas2NY1iysg6J9MzQSpQlFeG6x6vTGyjJRfoWAH0RtHguXs4YsE8dGlzwnvhBQw5oNmSVzptT
/QCkROvvAKwyCuILsNfHK4C+imgybmvhdjOcJOLBafW+Etg/n4OQG9JPxwiTBinjtWuGZHzVwNy/
ixvGdgxfUE36ExJdeLcjLbySEO/NSG5libXbwsv41vwGGfjso+ao91VXrGikSkcOhsEcDEuaRqKV
suKxlp/S7If3jVbDuqCTgR0bcrMXwehkTTkxmfyyF0esdhpjGOTAODd80/rdyaz3wyL0E2G60XBS
p/VZ3bUY69JnPHc4ZkgWn330CFl5JGS39gf97yul85lZMpWbrcss4SsVuyrMv+vYUFqb8MAhqipN
Je5C2zULdZA0M3YuJa2dbdLR/diCkK5fUJXL6gjNmKRQYG51lB7dpsGREie96nX1sPgB9DHQxAVC
k1Yfn3WTn03591p9iUrp4IHVZxnyng7Yrg2ansatINppnliKcJWigHLEEoEHt/RA7z3S2b0u9RQb
U7Z2qRm811NrGpHNiyxUgW3xth636chNbZz7SKDBhsIVAV/EhmpwYftCkzak1Mq+QldCJPAixd6G
UmemE4xJjDuuysyC0WJeP5RF5byVZHr2zUkLElLQpt0A6V4oE4Sih2dXz1sCMVmuaP+ZsIuYkPJs
FVn4m4DIfNgaGgVqUXs2edCh5cLC7E3KJhPMC0ZuCNziwfvYgdyT+kgS+QpolN/exMYvXmvxxODS
Cl2CKXJjIgo4asFxvpDx8bY4ODcLUGxU0P6CU7NOHDauaBL0hhl1W6M7a8pKL2E4Df+sWfvkAPFR
+sJwtPXXbS8qDCmbWKmWko1HGBj3UdATtf+9fAPwaeitNE2OfokmBsGIYm1IiH8Qceq4PI1r5BGS
nK+prRbkCDUMvzMLd60N0znaD8cfJzjCUHXSfHCa0plcC87oYfYD1O9XEdcW2mxZYTbiHkRS1tCv
PRgbiUrt2aShrhOf6iezJjxrmTJv7cBEgzhD9roRhX1cskWhkLSZdODa1aea4x+w80XEpSAh4t+4
bMw6LKlVieWUG7wHrL+On2oGBJT4hLfEfPcIyxNlVTB1HRcX1af/vDrECFBv0ns6tekyVMX1AjdV
PpKHTsBBe+kt8OnK2kMDWI9wlN7mtH9wSZDHMB/IdiAFH2zZ5DVEtde48tDvJO1o51auIRFSaVYO
LJH6jH6Wv7bo3m0G+SwbuL5XWAc2vZxLAuMowXkFc49SarSofJG4NaXm+dJsZD5bOmyWSDTxUZ9+
t/7fGjmsJw2QALIteY8h/PyiEwZ9Vn5CGJ30tn+ij8OVKeOhGx69nwJnsXA9ezcYWVE4C/bP/oo0
rTo5FqmacCyMsYuZV3SD43iUblcr1uA35z0qoUbkhiCq+ra062uyMLDDDKmA/wtFopNU1LldS9+s
MsbrJhstDwYH69Ni+o68BZz8zJ8cWp+OxGITvEIGgMPoiTwAY3/Niagwj2PCXphBXPKlJGD/101r
3Avgt3MpQltFwRicOfNICp+UgCTMY1UPGqML7dHSKzPU1Mqyd/eKQMvXRNJMi+pvgoigg1sUn6GP
WwJGvBVYnJnZxU99zc/Ezj4L/jvI7b2q7v1+W3Hka78jt637QkhrvncNqJCmYgv0gGaL5HpXdDAy
MToUIJWvwQtqsljiRKgSb1XXwevhLqlvwDBK+deP9dZxPV9zmxZ5O4Mkw5gsYMCno9tlGBm0BhA/
XmcOQd7sgvKIHXm1G4IwQBa/v3t0m2zidYbgB8WusQ4EEFQviTT7drgnGyGSpQ+6qAxdVp039ilr
9wJ3CJiUWXyE0Hcg3GHUzSogo05CdI9M+sHKBGTkhJm+7TbgusHJzc1+8i56jdWob937fwr9VNgG
iaEI4oqRQmA233o5AyRfkCyD+Wybtcb9bF2c4niCdLStvdc8rMdC4C9pq8QZhEeMJzmAoa4XyqJJ
8xoE5d931P8oCc3ouOIBfrtT+1p+gwLcWCI1PqqCcPhpQMR16z4+UjeOfneEcT0kJLeg70+nKERT
cb+2mL3LG2xe5vC2P9Om23BBVEZmZAEQENR01JUj7kPhKJgz2dnOQehUe3G3hSb4VwVnBKffEGvS
dcNej/LFEGxnhLJQ3O6gAr53dhHeDLPC0/OLWf/vtDsKhOHT9iaXcfKRTgkVnWo8kVlK5Sn2Tkk+
MOoi3sNIY9n9XV5BejMBoeQdeAWr6GWpK7GGb/8L0yUE6jv0MztrNZ+FfvFRy0xgZCfDQC29f5ZO
pHlDLwpNqbEeFTJOFOqzyUvRq8dOctiCyTcAXNmBnSGgWzuDamUJEvsB3ZleHNnrHsiHeG3F0nf5
oiF1ha5nMClpFHOtlcgJtPVOkWOKFbB8kVsLcCggSssO6LIbjfyp/5pvgBLZ1NeEtcJ+Lq+jX/IB
apoeGJo57IAfDNLFAHDLZqvHwIt/Gtn+M5Pk7jPNUC6u4zpic7QpfZBWF07mNPlnb66zDhhDgij8
mAU5hUDdDgXy42Hl93l3vTrk5+e4vL/CXqPhL7dbfuIGVUKLHiaXBKsx7Y3fFHDLx9DhNaWBVmFu
zFq93TVSArzZ5i19ppx+vxdZi4jnTFnVA2VpD/OESxAnJux2qFkejcybtTdQpZ4butocpRUpRuCp
GLlZxnc53n910adON/33iBGLlx8uCXR9tMEVcJtRv0STdTH4USeOmhW7Rf040+zV6ed95HdAs70W
9KMHWbYgI/TXf6CClUlLyDmH/TV1eO4yXwoIcZt+sZzG+EHgst7D41Ak6OMIlis57VwJ7jMvszJZ
ScH8GfzzNr8mAjWIPvE+YaUzS6SqzTwZSZvNw5zuch52/jJr8d5kYnuC4/QFW9q4PliEyrJgDTLf
EOiotbzhqaZpRaHrTJhLBR14uv0APkJW0EIGD0x9ZAOqCaV+2XIK36yF5/R8nThE9pEgU3Dbaw1+
ewasi/znG0bB70PM7s8AisXYAwGkVhIJMkVBFgla2eSESzYChU9MlVUxaSzXVz3uvjSjPYyraP9H
/mFyPoIz4OBUX69PbFXxYbkFxnmNSW2qf6EyWh7QfE4KhJAtpHoubp7PalefObiH/M6XBLx8qekE
5Iv+vbvuVx3m36kJGoxjQ+9FeZpnMqca8uc9uku+ftFGWzJqw3T3u/9Tm6oE3pgrhBo5+havDtiI
LloCaOmUgEwXnAF75qMJ5KabnimyBZ0hCZU+jXzxQ/DodapwIcPo2WJdVFcoHsErTHdYPWFJySTU
bZiC8WBRoVgNkZjddon11ASQP9a1bU5qzJMzFJGGnHpL5+nIR1sUgWzjlt8bc+o6VJykeQxkhto9
ZMa7MJ3Sy/nsHPMTP1DzV49+u/0GgO97fFOELAwoHLhWL70365dg7gDXxBMlHbwKGPNnunVeFy/1
aTwj3QSnkkl8+Sd8bMa9gHidUSHkTQkLnOcS0h7i/dH7lV71GQwUQGNKDGhuu67GrOxkmRfVjTEt
2ce1qV44iTKPTafnd+vqE6wUM/tSOUSGtkgPsrqcU8E1UuDksVEKAIjbDcyNkp+eSvjN5/Eh8D3s
MEzmoH6NJYc9aJZRJNhuukQFk2e7b0nukM2pZLKwO1URbAxksp2t2oHEPJu9PhBpQGSpHbeQzhEo
QsiLfGkIwUqMNPVUrIT11zlKGj2cMROaJZYsfejWOSbV97VtnH6rbuyax6TBUfz6kEN3EuG3lcMI
oujikvfhutWgR1GrhVktNIlkHuinxTjsW5c6InZZOUwMVhXdi4joOQr+o5jHUskQ3a5hPhrlTVVG
UDjJQIBYa5MphBZ57KmEaxLrQQY36hYw946NgQ4Pmy48vJfLD/LV8EgJv3lWF2VRmYaax6/HAYo4
fBciNjf6mPOeiNZMSJx7nDNZ6xmt3wG2qBdnt4kVXU8RPNDAO6YHqagYmwJC2XSxkrpDp/x8LFmi
B+2hvrOZRIQqr0O0AjKaXxuGe7hqw5SNS/QG5AyfLZvjW//jWzkQXYRMrSj5QRX+nG6rof8+zon6
f/u2/qbsi1WEUQ8Wa07sTkPndXYo/mKQijXj5XDDbbnzBjPCJPqc0POk5ueBrSzIImONgz+GLwfK
XHj6uTD3XRRz4uGobQ7AxvdEM8YdhWgC562m6jmXiSxQFnBYkBz5MPeHKWP3Eqn0BKaXby6+EgWk
BDPK3L0qiYlnPuBVN/y1Bo54JmnTSepLia46d/g3fT8+UahivWIVybDDRZExCthwijY4WS302B9f
turG14IpgrN5a9lXSpMvvT/dEgTF/HiFGgS9uUz9bp2TTCh9eleimR7erV3tYarCeBI2Uw0pNlCV
V5xqLP4SljQk0sBmrEutEahymPswIjRocQuy3+dYmzDqFrsQ7KOYD3BqrvK0DoP8K1Vv+SSxPwXD
3WXfHINWvdRBQtD4r3LZg/2HVdDpYv4mHZ8ZPLDif6z3hsmh5VTz8j8Dkvxbrsdu2lnRKBF+m7M5
PldCqVLlXs7vljmUjKsuC4f1n9BQmvBbUYA9TpFe4W6iFFvbi6aJWvUkRfHdFGtCW/5tV2wnnCjQ
Y1Fx8OWCbfKgWB2a0aUoroBLWCmAJOLP0TFz9FI8DNn5pr5vGmJnFyd5frTwifhyytZsOdsAuSHg
Sdf3kcm0AFAfY4tbE/sErmN5bSmMRsK22bDe5Bo4HuCJo7wCwtDz/RlODOkKh0Et3fEJ9gcRbWPX
P5FeB9qBOuVnSCSJ4M6IiPeW3VbaDDp0dNcX+hiSF5p6ASDv5iVcjkZJkw/qaV2yPAWFRQsFTQs+
DcS+1EmCFDEGj8xcVCBPds+nvMzJX0kGl36YAQTZY8CDVUGH+T4PFiUeP3uPmKK82aZLrRMHIhlz
wj79tEYGMFyfuctIF8CyxGoncVnIvnNFY8UsxItks1qeV8lFl7MmMCKbS3N4d4RRX0GUxpLdzrXV
JBPhbWUjpV6RkfgomA04kgXTkSJeFaDrbyQaXrIFRHvrSTLlAMLWd052ZW1VRa5O/4u+DaY8Kq0N
zP+6CQv3P0vAXjToEOCd9feqjg60RN7QiZjtGXednJ1VkrToYKl2Vb2V71iKn4zJTjigw1+0X10D
dYAWKhTLhQgye10/VOD7zPGjrvoIQLIGklAUpCOfefSerbGmgQV3g4at57Pw+/80/2jbSO+J4BWu
EwJkSb3xrP+HzMn9iV7dGMKZFI6Kic7d+ARRQFjLddRIfhX0wTVy6tfT+86nVyTIm2EyvP0mzfSx
DxihulrUoTZlAE7gJA9hFmrAYtgCzwpFyincvD68swGcK2NViv7wTHU/OeKzp5YCYfy69zgy0loq
ToRNM5e1hOxEq4nwWWBvdnaqXRR7yLCsDtl+DKSIiwqll3Vlgw6/OOCQbtPZ677Lvt8ksOBziefv
fFjsWvhWZxH7j/eWGdMmf9bHYLj+lyYZPOrOyi3QU73R94IYOnXuRtju0qCx/aQUV63rspp3XDaJ
MvDuXTkuYUCRwvgLLLl+oaLj+gLaXbumrkbyTIrwpGfLVLCB/ez4aOkjk8n2YrZ/p8zkt5IGWO2T
jv3yf+a9zl/JQgV7TsD55NPZVYUGG6mBGkDtObDO+sY0xkdrPlZJIj98HYEjwV0N0GjysFbOyBze
ZlF9tzEnKhcCVYJx6oof9y5cIQzePf7RAAXIewu6lXrZsoaaroJWLwwHi+4YS+5VV4kquZQ4RNvP
HTwhAPss2f0yPlwT2TV/7y+sbrI4ywDaDfFJW3kSm9qSMFA98jGNEytsU93VVwkHLe1mo/MffUlV
Hp1n9q1bjXbjmnft1Y6Ty7Uik3dD63mNAL6KMq6Ezy1sIzu5MhUDeSBYjrhcrgMEXHOu1pAhRhGS
7We9PWA7DxBTAXt82U96lp1Z9jjo6vm/7mrfE6u/REWQZQ7L0bHn/2VEsFNX++KRm7/kCNGNZcFo
3WkTHfyxVTx+T/6dZrgJaXaijL0v3C7ylaLIYJLzfY0LJGeDeooiiH4G+EkEY0J75YdH8bEzkpv7
mDAevDuf9rU17EhnxQoxTQjE2uqG0B9CIRV1Qd2kxsvWelP+aOUMniffP3/6zsB4nIgJZ0yYEb/J
vAD21yOjhkBQOex7x0c3IqREGCliFzw0l78NdaCGE4S4/v3YJPJmkU0T2613AyDdT7I8VJlTZRSj
V0xt8rfHW2+xXewFnYXd+bgWA54NblCCvnsIZHnez4ICTkJrH7NYgMVwjDdJmpFk10vQdiPVI8jA
xgIpOvpH/KmifyuWPzIIQlqpbL8fZPhYSu0IITvX7UI/6uJTg3FSCYVU69nGmEawliqVAFpqwqHp
qr53PP30AGenwU4Q+Ym6dCmbpHunc6bDduCfmDR/ihSVqZzR1e3XpiztsD8nFToZEnuGW8grnsM3
xqZpcClm3rHfIz63IRgBVWPQkYNZUhNQ24RLwbG+iihDGcIFAeMHBCXQo4M3yAqpuw2cd5J0sa22
9WLg6Vm7bipIYKERcw0h0FCQiSRpJ/E+xU0sX7WK90/qrH1GsXuBlBbVDDjFjtNBk47Iw2qsI7wc
Ww05O2Pb1pGtKPzT46zriF+DkR0KzVEOKEBA1cc0cba69RIOgtvVo61ArRycnXCL9ENFpTCsKcng
JgKepwQU0KtRk555b7gqRxYXvsrIfJi4joKTl4w1gz9FOPJnXcyQQN4kBmwROwyHbs9JIkdDi/xX
rXOo3OQbZ1Tti6SmlaEo+URzbykluT1/JJll7Xk3TE00xUTVChT9YaEFEwhrZxOGJD3cDHRIm9qd
L16DYjgPPnSGb4YYtoF7+IwZtVl9iRMLDbHoaOWd/OST7kCw3YB2tzhCtfU5c38SR+cmXAn6BVvC
wg9msgzLdMBXmXVEmGuNe/c0LYS4bZd7EB4QdDUg7qsk15qkvbqyi9kQVwFHqT+OWUUPYMmiCKGr
E4uDG+qRAuF3PEqN97ZrOpL/RmsRbOPVHmQRgzzTbVu6JHcrxLCf7m4cbswj0CSbOefvqHVj/+PK
lw+h8jNjzfAMZpD09afTZ4PxJJRnWtdT0p8hRYL16ULdLcd1g31HeMOMlxbfWYp37p695a46GVxP
0TzFlleLu8O1w+c7daejwE3XjsI6T8iLA5FtkTIGC1xgmNDkhPaD4296b0Chf3d1onmDyqGX9Nbb
A3KLw67wDd+19LV6hEEWA18j9/jmRqgciy0g+dEcwJa8b5em3C1qFxbSkwBXTWlBrHiCBnLuTEwT
BErnOdflKbo26RXwrbjJTAnvjHo4gpDxVn0kaDkoDoWh6oXTRnmfjKZAmLQaoAZAlom5xSHBsa5u
VKj0kUOcN3EPGkJKUKnFQR5ev9Laoo36kiYjfsptM2r7hyq+ByttX7J7UiyDPJzE9UUkF4e6/KI/
yUZS2VFWAjQSy7cdR8UJh8ode8hf7iZugRCa70utB6GHau8nFFG1xG5hSHwJ19Ig9YVVjPil00YD
EbHy/trAo+/cxbMfoE5S18WKGLjbsNJUanlld3kYO+5MrHxRpenZPjQk0TRCIzzwXPP/f45OK6Dm
3hMFObNcMoMn18jV+lsi2CVjxDRNGTElbzqAv/bU4vnB1NYa+IdEjhxG9RE4fvhv1xh4FGOUa8zj
gz0HYjR35kVToYzuo7vqq5cZfdPE4agw53Q98zPD6fCofyXJ0yCrhzgtC7E7s090DmSw2U9o90DK
5Qm0vTdyeFE3DH1Me1PiB7/03AORUmzyzplHWFASWf03aB3JRD1Kq5Y0DA0OOfvhQAoHkTW2q7hF
lCu6nTNoqXvlb7Ne7LTbQRRPHTb0cXZKXcrP8OabrVmZjRcSBZHmBEopfoDtOhf+3ezFhhlyl9uR
KKH4/fHVFkrbmtWWfI+YclJ3g61pPGEvZTbVHMA9dYtIAggRSZOUbLmZML0MFHNb1Y9NTeh/+4NW
tDAuPH0SWFBb46u5Z28KRKH5A4n4Ryw2NI0gAEzplpIGPgLfr/GtUDkK4MvAbMuJNRzAm4YQ45D/
t83pgc33w+Hci7CqjhhOuUfqESLzxc51FP/gZ53m1EzzcUDZiG4nNiF2KbVN6X6+KSnm48rC8Jug
2dmLxqEig9LdbeBCiXu2ZxIAnip1TAzI7SFmGXFdxsDiH6oYzWB3g9umeIo7+kxZYpwRMfhuiYXd
7ByP5aivvfAEEq83bvA4lcm4qELGJWsBLWMLOqNsbzj/U0gzD2XUnSisjz/f/ZrMHH9uFMWoLZcA
5OOFp4lhYOxUzArV81WiH/4NItHSYGafBi4U9gghmXgCe4dK5L5llCoqwqOEogz/1H6WlBQF1CQX
A47sk9CzIQQZPS0TOhDhQkqf+XliYCdkSST4q1Ck5/ORegsXsCOhgk7MELDdGWZZgTQhppmMyssX
Dq5UfSd5aBdQSx8H/YHqnP79KEOzcZ0ApcOOBFho4gbwvrJDzgtlM7jjdnbp/NXDju8u46sKFGZl
rJYsfbTLYAc5nzMfgVl905Zfv7LOxZVcIOAVOuD+/dqjGi2NbLY+1B9E+PUCq4YtOARyiOl434Fo
h0pVBEmMzuMbUOzVN+dcQICMfDTHroc2GRvFMB3l/O75htPXllEG1f6VEHNXhHgbn2gelZdNIvTe
tvFrTAvXMFWVfmZoNxVcCHf5suxAznAIgQH/+UaEm4UdoeXyuDD4OLRtvPtqUHQzFYHj4vgdE3Fw
0zGpzu/938h+4sn/1dXlDIVebKlOCXEEcwC0iN0uhM6q9B+kmHDccn4Mk/21JrRfFUFqzgiuNoXS
IpdZN13z7EBfgneswCAjcd3MBwuRjB8QqXehTmgTq7Tv3KZyikg1tImb59GpmpyWDjAhD1QzIoXR
HRa81Q8+UZqiWMGSb4yANkVXXUUzRObKkJmPjYt6lCXSkWHA0emqtL1rlPLY4Cn1z53x2umzsNCy
rfg4AKkRVwTbndWEvZ791CgCses1MZvRNlpP6V67gx2Y14VlZfdSt6SD63f7ivgKCqNchpXa2WLp
5ccVC5IuczrMahjPMPlKHkSb/kukV4XjBdiZ0XbWeNLNUNYN3jpBuQ1J+3PafR+aysFT/4MhTeN2
sNq2/34iSQkUfejzbnUIww/Hk1CuWJ+Sk2RU3HuRlMduaQn4Ni4gFOkpL4fH0qREduGrP4+vxcbT
BxkvHMQ1l6noeApD+BCFoXSUhWwospGhF/e5fbXSCaf9J+nTYfp+vGrexfFAenuh0HDwp/zjv2re
sWH8a8EjLK/94XegumBjVovAyfmfe2BT3i48CYdQtzdlnrTtcvYuWkAwrvkJfxJ3/il2XzBpMq3S
as7Gob6l0WcbZZ50gdqANY8AAU+pa+WamLClSRdHbFbzY2DxdmBDbN86EO4NfdAGmlk1yabSMgHt
X1tcgI3svpQycBXJgvTpAZrVVXBw0qTDCsLhFbRowmiKIb8EdXyagapw91q9fMOlIPGc58etNfbB
rcWEGJ09CRYBc0k0WB8uvCC47jnv/y3fQSR5Aji4ihEdYEF7IEiPotfbpVMEtW5IO+4clZpnihRD
u0OMgwrHbEq7UPeSyW65H4+DTrjh+kaP9e+4xtGPicCGZP5Wlbojgps9bJSYIMkfKNBPhSmD6HXQ
M0LO3p1fXTWbcM9Xspv+OAvCtkph8jpcVpAjvR1nr0L+sd5nHIj3KTpONuYwkm8+IfSwy+N+4DOx
cM25udcLXznWWEG6unAh9STyTLps6+SlaSpW5XBRbX7iQsQdmOGqVYy/P4FPW4c2RA1Q9hpf4Adw
8GmHHbjMrZtOnI81B1hC3vyZvmGfS1Lsf/AcreNvBcR73bDBugel3DKmWCFgOGpHNqfI+aPJJ8T1
tlZMrijqqLaU1vXNbtXGhOkxWAkdxXerI9JfkodypznTEk5eDox8tKNWiDPabjYZ6MLSmPiS+3nL
H1gUzhj0xjNuyz3w+IlJJFWzxGSw/CvWau/gUGk85amgq3ZAK2yk1eUV0OxW50bLX6h2c88Ua6my
UODsLDPuwAoZuLf1Lior1qbg5R0XP/2FPpnTYaw55Cqf8bFhmM+Syxl+Ug4B3MbntCDEGGKrW+XD
hOd4ito3JXPDTE9VRA1gE9Npk2X/eWgSC8/QOsLjlzGyTDdTw2YHxadIrjsUmwtStFGTJtDbVme8
+RsSUiu1PE67wZCbErUZIS+xtk6mHnPgkiosqbDbD1H0HNSEAffoBNkp0ZcgCbt+YVlfgL0oyYrY
tS7D8VbxO+OC/tkr6eyXD706Y7Til1mANE8IH9rJdTKiw93eVskG/T6/BlSygTG/5NiTbyIl8FjG
KIg3aw6+uelZZrkfpLc2dnDqdW8/efeawp6kMPEpj7wcRb8ZH3EqYkzQN0Q2xfKR6Jjm3eR0VO6j
SS67UYSBIR7TLW4aygqk1Bm6yQpV7Vx0bLsqYqz24bZqVScgtCURm9X+Vr7gZo729/EfV+k3uGv4
mVFrl1e4LBB12620fHePZK5tGGFamKCLhdCAJn0iPqxn85P4A6nCocJ6esp5des9VL2Jwdo0Gaof
obj4//6kgTAdQaPsoCTnqaITftT2OMuFDBZkAxtGRJjp8VCVUKavhkk0Nb4InGm3gPJJI8afQarI
fSXR33vLlxQQtPxoxRj+K1erQkSVO+dQT1ACQyT0ZsiZtzzvRZvS5ClcThoRojgptDXs2myX64P/
dgw9HcsO3nAvrZnqrqZabC2SFb01FAuOPzakP8RaOjSzNxW/dE0GhxxR/D/HI6DCMxBnLN2A4m4b
QNQxAImHpzQ3pUhcA8lGAGRY9roVyMUwH8GQe7TjfzAkZtADWgZju1fqa3gfasODBVyaGuWB8KIa
tTaukQt0rWe71nmCoKsbVhghbmXpXDpu/Uu8nwFt5cPfisdCrfyzL50Hao/6Y97U9Wbmf4d2C/YY
isGPOONT4tITYhByMAkqrgv3tqecT5L8SxE3OaWQozSoa486+fAMJn0o93zmF3LIvBvOBOBO5yfb
4xWbJFTSJ7HqjxE4I+CVl6MGXNE6kSrVZ8n1c3njUY3aVZU/hPUAvhW1pUqN5ntgYoXgKvyjia5t
1kdDSbTLmcH2IYWao4tMNZVmrPy0KP77hOezk/VxA0CWgYcyprq70A8/t/CzoqGq5OWZC21lhmeI
lfycQ/WnDe1zs3UKA2Sg948RGK4h0gwGnapzmqjiETJTgvijJ/YiKQJfaiZzbQ4jyE4gYmJ4KemF
hXcbiqRwOoYaLjxIYFP90sgmMI0xfu4v9acnGKEQ3t+sHsbS6nhG6+in+/+HEKMZP7Pr35Jt3Cef
hQYj3862X4RVjfDErmqq0hlZtJlGFIhwgLs6/7hXiuosXpVY7BL9gLn467k1WBfrLqrGQlhC+9CD
1YlIFdqv+bcv0NRs569O7T0uURjgIme6UXlvHqc5H1e3B2gTjhb9OjQc9UdApEPpzRMW+z93w4V8
iR5SlLB5WwxTUlRU4NzmUWWcE8rzKWVgVRB/Y/YBPqelTJYmKhdH+i+kvX0bI+q9KKsYatxT5Brs
SWM5Z/hEOT5ykZ+WZsJ0o9RUe2frp2srC9jFqqQ2vMjB+mdXYqWkFPhvSg75BmZuPNUyp9W+mkI4
DjXTtS5biDIfrdOU6ZCqoqfm3P2CO3+arqr6xDJ7rZVqQXQpkEcFTY8RNPtigK3viZ0GS5WgaMWq
3Hgf2PfLU8rdkl1N2PVggj592DlUjHuLNkbhl7d/u+4tpSfux7ZoL4NiLb3PNP5ogvhkmrIOZclR
gPsnAd6bIvmAUVjL21Uf2K7d3PIe3X6+mbZ0Ltl1skeQuWZKdrX20xpnSsgbvyChENTtJbFM74/k
CTKG7LQ2zzsjVKR/pvloIpwRdytquouqnBmQqakGJH0X0oZceXvaflznjf3oc5BzMITubPDtDCGf
uM7kMJ9PbpI6rj6rSLjJW3mexPhu4JJ4tcP51z5g8D1ApvIRJnYwOV7RzeZ0zNcXLS35U67lSpa3
GsNMNgfY3du60LUfwZZEJW3FvBsTbC8x4n5eViwBPpfSx3BuFEYuAHpgYXH19o2dm/TYyZB5e9YW
2HPB8oiekFy1Wnru58hA/GHmoHEvTtEKzV1prG5WvXRhwYCflUGuP4kKorLjFwmolakQGUIqfH3i
DxN8pTKguLpth+pO/qPrtlWD9kmFM7I3ECxL7UeQh/E1d1yNIUfiswiKYX4DAOFl+SjEMiTXOeI8
UDYl/cjZPDP5RGyctWx9a6w+BOyAOooz9RyAY2YeDCza1Awu+PMFJhMl2ZPsEz/ZBkItWYucExO1
lZMl1fLEH3rcc/9U/BNBFTymWDrn+ZBciyx6de2auJGKOv4H6YZG4LU4S14u10D1NoEHlBx4BqtC
31qxJN3p7kJ3s+DqTbCS4FZXmBeLyKT92V6hD9q197GCVvEjl8nKwLbAS8I8HsKhnRmyU9vzBFbL
Sz7627SIwQGR2OumINfE511J2pG1KzQJ06KUT560vbUPK6dEez6f+zyabpCEg0ebh0ZxhQDg3uTO
WRW3i2XcF0+2aTqajjONDYUf0YF7UN+aDdfm8JMgcvJQw8S3Nbip8tQqVOPJek5ZqpqaObP+lVgM
mORtnaDCRiCQVacVUyW3pYYd1avwAYstRnDI00UCMw0qL/CjXV9jIudrYVFopZyl8fO6c0ilSjBe
YkKFvp5/VNuPvUVMluXmXVzJL8xxHQE/z9+8pRlVbBG2yYqL0eYfBB96WNAV8TzP3/L/F7qc2ZWo
brpPrjSRkpMxARvXMw0PEY6o/s6Gm+5/MOxw93yRFhJ3qQjQnLOvymj/Hu28jRS6Ok5CcTWFIlG1
u9oldIQTpvEdsBaC682NrlhULxX2QcmP0WnZIHHzp/MSHr2go7QPJFYJRwFBCpsErhMo13afTSyM
/VgUtBald5Xo0zMXaKbAnqW6mWykK4/wRm4vYEWMIm31k6w4ViinaieCcURNNd38QObqf7xJdt+C
IUySLtThWeqZm8lfcUBx/xodF8SrUxdn4X97/QAUY/GQTGzvlf5xYxMYnnHorgBY6OLwTzung8v1
RxtACUui9J2g/ydnBOuP52dfpnFNUIbwciBAd4cXqvJ/uAkIR7I52ib/4f2TA5TebRKWe5ACbXEm
ucOvuipWjPNfcTO4IYfQXiZezd2BMCSVjO7PuvRyH3rUe/bgH89ZwqqIKm2c+IjVHSgAhzuDw7II
vboZAZZ62na4pC4rbxVlJBB+fstAJetzAa7DxfqjT3Q0PqJg9M1BI933kFUqgZ4S1Ff0ZZKzjNld
kwQ/+bG1Q1pfQ+5lgUeeLrwANUOyprLJuCvvtTtKOhUg1nGEo71ianjr+CvwrYAt5TKMJn774b0c
y/7JCfiFm45cw+PYZwk+0oZSJeXiklN0eAiJuGINvLeDR7bGW/ZaXbGAb24nkCdNBV9QxPntDI9W
oc3RUjnclP9RldY8BzB6bcugg9/gUjcHj4ceQPhRzcfKrrR+IzPCfqfgf8J990VoeanpGDMMBTuh
+k0AUjSeu0DvDrF9NEGI1MJY1+c513zLL739gbReKY+RjSTcFGun4BUkAFCP+z6l/XCRLMBa8gfG
Wy/n6lq3HSqXhBtcVZoAp6HSkQkJB94CvOiDBHfXRviH1p6VSQ+8D8WAblB5exPMFmi0/a9n6+pP
jlbpfzJ71dLEOXKKxL/L/y9fwURNkY0pDhX+eXDmawBxC4EaTO7qcd4HEjHR45dLf2oq/dlmw+Fs
cN+YO+wMH/+4tKLatjdDC/sHx+GFe9ZmNuMy5H8BU/t5zXoF7mq3xquDIvoVkj8oUeyyvYHY+8oX
XbD9kYlAmy9x+HOKnNcem1Cdjzgy7FI695GdSWF2hmnhVvpFbB15smib/81qrQX5rg4CZ6hLqu9Z
bvpqgNuWnuo44Ju+YdGKzECGDg57WgAwVAJ0TlvreCGIlWxmK04tmzgs7q5Wztv6HRuwJp7+LBN1
7b6/sdyVYw5g0+s/kWhh1EH49PttWANdsU1KQUJOd9e1N5gYnfPziV8aH2on90VLR+iY61usCLhV
OED4pDGLndOs4HyRAacCp7NBlE4fcc65G4+8S0czsvMG9cYpt9ziolRfT4Ou/M0367qGyhxMfL49
1+JRLjEQ/AtqjtQluwor1RfluoKOnWDpfFgx0wZjnPYlpz3kDC45bOc/ZI5GonWtpideSNJvZXcd
/EH6TO9DJWece8uJqYZytzF4ezEtxqAKl9JMj5hUohnGIsFD95xJPuFMdmkoSD+tWCDfdEKMC+qu
1Ucsm5DSfLh/505ZikYEHKUWpoEK0rGLGz2Evm/Pb2GtyKR+WlHT12N8sKzMAaa16dJR5pVE32Ld
wZYlJ+4xR/pojznWYxqy+9dkGhvtnmhBOwPbL9AdhuofldnNUX4nAzE31WPc7ZG5fbQOobvFYocf
gX+OkBGS9qRVbTmw4ZmFVmvYEltxxVfkijaQlNh9DA3Q0tHzeIbqz+DGoNxYjfSrfnWhGSFW8/Cj
VwtUMq1y0351BTu3JV8qTzec08/eJ1g7dDDKV45Y2N3szu0oz3BFSi9cKqm5fAg3DBEESROtoWpK
mAMU+Ewt/Dj3AsM8abM6t5no0mwXY/jmpukyAStVTvhe610+QAv+X9kFpWay3052FKrgbklt+6iz
fiHb3k/srfuaGqZ6dJW112YvPTLF9OUjfZdL2Q8Q8HmD6JY6FrqFix5unL2s/pfQxCU8dC1T1bxz
/ns7B4qVtSQ8P+PeGv5JC6LI50H7Oc8HBN4ehFrIlVngCiPQqQIogxJ9i+4njh8Z/DG5CxDz1XD2
Hu/5uecKg4UACR2eUgtkjZexDiPBI60Fdl1EYnJ/LW5O40kwOnnKVjTPFq8FT7LCSEjo9ruiPc+Y
QeOreUuN41uCIpK+pFdyx2iXfB9uO+lqaK/FHjhGTYP+CzAz6FBuho117EKnjdNsr0SQcahS+bDf
jGBKp9XLdXNSfYHBE08lCm0cPHMmKf38gG+IKu/czF6LDxk4uqjNQ/yZWhQm1QUCnepQjySaroFh
QkcqFYD1ATYMS8jZkQFzoidq2Lw4X3ldCvjUGDHlasCHnVd95uEgEZWwMkNCw6kct1K+IWnjSao/
GFtng+goTi0oJtkk98aexYgcYKxdfeW2iTni+qPZKIB0RZ6FZ4pbIYQBU1evYDMa5EV9cI9qhKlY
QD3PBxT0B09BQ2BlIrvfCGx/Rke1JDNvcmIIAQjoSx/wKvOI6BGX09RwVawiuWkrv+ZOZRVg+Uhh
KcGNLEqyeZUyx1hIFjcYihrLjGfBI+AKVIbEIll7HMobAB/xz+PPniWI0s5CmdtB/1dEsIWklVgw
VvadswVUQ3d3LFcjgba5u7ElltuDChbkxQxRyjZEouFZS8EcLv882Dweu8W+toXq2j01LFCo4bK3
FrCyT4nAf/fkxhwowo2Ou7BxoSk0q6D3ndCbID24WWqJjDFHsNkmIfSnJ/Ad96E6mBIdhFb9ve4M
t+QSKIrI1JuLed20lClC/stwVuULh3Mc1ToAgQXSuHdd7SqK6ZPnH+19LS3a+ik2vvcgyVyq7n3m
v4RNRyQeYAIoSdxJAig5YSqMGt+jAVEImNodH3XsN52gwelSMCkr7aTf26kyR/T0j+4V8Ee/tNBn
4OQag4Sz2gwfJwkgB25kO8sqxD3/S/5fzlEUhto+5Jza1lJEOrOlqkmc3jTRbSe6mEkikRIl29gt
xVvdpaBe85R94O6y8IF1gXndK/Ak6u+13kLnGRKZdpayt641f1Bhwt6AT/DRKK6F/eSII8vn5Sku
jJAUXyLtybdoQLqfF+Z9qjIrxWZZ3KCNxg7HNFGzuxYhK/tixGt3Zq5p+w3l7wORyBrs25+Ha+kC
tbOEaJXL2s1Dd2M+QS0mknJzByqyE5bDsM3gBqv5h0+n99PhT5SfkBK9hFoyJ/Z7SxXlEFyOXmsb
86v99W16AWFTKFHO+ntoF/cHkBRHh6Tr2KPwHMWAIDNekkC448E91XR72WXLObOg8a5yr3pBU+MZ
f+BSRfQIbkk9p4YYxv94E+cUBwxCB0POVf4Tmw1i850b2UmmswIhV0sT00NHilLwUVw3IehXHjmi
8OUauq12zjgiV47oXWtribXXYMFXw3sNfQyzAwKcCEAGCL7zN10EGYhf2v49nu7By9sAF6Vs+n+i
0YQNGioIKGLsYNnZrKwSmJFQUV00Qr4cgtY6BArSbe6elDFzoXdoKktIbWvKyQjgoiEnSoFzxfvC
KESYHs5xgtU+MgARZg0iA7h3O0gvYwiWSxK8grbtdjDLr3jaslxhdVilMGY0wUmMOBVdOThpOpau
s4yjIPDOP9U/WZ6CfzR/hPzD8oAMk0sEWjhv0b3wM0s1+ZQuE6ChbxCYH0VdWB2p+o/GdHdWXEA0
9s2gdfzSa//rWYg724J3TgOpEo8BtyvlAw1C/TbJut9Zji5y5fxRXJHMt7Lx8TRMfhXjlWfWM0DJ
4w/HzNHl95cej4EvSmI7+eIqrVnEfv/Xi/G69Yf5U039hjN+vbzm+VvkqWeGgUATKf4kKmZYkRXB
OAnL6BrGDWNpJnFtfdv+Ne+wAVPvxPpWhbyaf5fBOMyuOQOF8cN7KLv39svM95HZgfClXtpqaYy/
6KyOup4mcrJflGLFRI07TKfGspch0HfPls3dVUBMeG8aM4FqaEZqDjmVJTNlEtcuWjpLNs8aSl5t
8+Kf/BSaOesw1j3Pl0uaMQmTqvjUmCSKkX1fAfVFmU4dJ9Un/Az4mCqa/UU6VODfbCxXorQ6jkYZ
SjrmsdhX1JU+kJvPllyiMhOe7iEpPV/9SKBtcMR+gqCzy32Zqkc7W/1KtZElWddhdy57mrTzLIl9
60Ynih4ngcer4ui15gEi5T/RydZX+idjFiyJnLChPUCpCNmoIxkAcDM9OM3qq3rz06fGAHjsSXmw
gwoagQ7MaGdilO/tuNtxul0x8a04XBI7Q/Y0EUuFJEH/ZTI41oiiNN43XNhHjuNcJT/ao03FUqUE
J77jrEq6c5ml9nQHC8wwSpxF5OeTQVEyhedQ/xFGZPRX0R1akleBUYYQYQyvV9X+4wu91Um5968E
FXJSWJfhh+YDbvlYQPXZgP5zrM0mEZBimSKVRPWVhe/aT60QnUgKszsLl61Jk6tskE+nZAMd9JzV
GGR8UHz8/fpUQ46QRMarQ8osjqGqT88zwH1tnqF5Cn/5Vw9aSMM65UsWPUh70IUm2R8zVLd9xQgF
O/t2+gb0gMTGyb4K6jg04eaXS/d5T7KDHQvCnDbLSVsyUox1yaSXo74PIAkV7UEgIBcjdxhus261
Y1ZKu5F7pUjD3QJlhNhmarA+429OVi8NbxwxQp7L9ON1zuWrhVBFEl8IIG4dPk1Fp42kmoT/5jm5
LyL4ovSvyJ9po7uy1Oe/MtQSrvLQGZ9aM3lTdH+vI9kugvtYc+q8rlhp45/uGGt4DtaruaKu21Jz
gsd1MYNLbHnEh6fxu1dLMUyqCUnEsmht7wsf6/LeH6nLG+2SWJuOtSM/WaPEmxQyakhjB6YA3FMa
i6bmIPLMtliVFBEla9VqMnijfUwLcey0ymJRaZxl4GSDjF9du0QOP+RhQkHjdn2nL1IqIXk4rhT9
MPi9L4QqR/rDJTZkrUBJJF/KwhWdAoCzWfUXtxGAKj+dgznCtDfWfeqtrmbJoGO0Ud0z2a6eLkwQ
5bTX6ovm0q1GmyOfhLsoN/l0/8D71n1Qv7nG/lXsmAiululjcK8jTHuPXQVsNy0SOb8C/TOT6M2C
B/wPOtrhogKJJxbOJdgGc4jz7ZwK9S7EmPK70wAQKWL7LEzB3m242rVe9Oln7oKNo7Q57gIchq2f
tGC4rD6KwJvM1pXh4BZpsoaZdrOiSbMPO/4g0n0dFRjS0cqFIGEaGxLUzdexuuxLpIULQHUncXJb
KRO3SKhDqUZdDodCOdGATusMdGnLu4zFHRWC/G6vOrvS4qvY0/jXdtpIEko2gIBSRlOCDedWlxkZ
vxHehkVO55oONc4q7P3mfL8wmh3qQC7ScKHDVq1mh655rEg8vWEe5+uloN1I1pSfEKtk4EdaCEe4
wmInD7ogA+jMtk9rGNPH6bEPNvqc9y+iqwHTU3iG2V+dHEPh4ZkVogqA3MS4XYWBiprytd3SiqGV
juSuoG2NS+JCuez+oUUHlLbO3IC2lbV9MoSISmxYWUCf5g79Fd6X+kiSEIDfB4VZOd4LUg6qQ/4U
pdp0KTCsJV1yeNe7sCNRpg+h+8xgYqzjUOGw+jJEy3UfjdxSnyhaYJ6HO1lnFmcN5p8CGUDTRsYU
GdAd5F4RHS6zTboNkAN4HCXiUMMLvoIKKXTq0562kTznAN28qrt5XnawRkBbbifiGm/GD9PQ0Adj
tunsyp4o0gjBh3lhN7IgmKTUOoON//JLcoCU6Rm/Bbr/Tlx7EwAG45Paz04EB4j+WHQI26rHx101
BblLOul2nQ8i+kXJjONdgY3IkRppyQVz0k1Da+eHpUrdImVtRzTzvJTFiy8nP3xQ8Kj/ko/ANDaJ
dvutLAKX6GcscSYU/mXk4LjJHmUKJjsqKJtPL0qJXxGVPdDV+aYaefxShfN/DUAY2ZEr6ZQGoOiF
rMS1VZjB2p+dL3GyvXnSrjH4F5WZXrxPElgO746KQqx+XYrk3cJZ4uzOg/R7bI0veR5xwBJCsqkz
NeaftyTb/njPf+4Qg9KqpbMicGFNC9+m7qmXazV+34XpRsgLWe5hucrS+gH2eWtnYB+9CQyuP5B3
4qK+wQ+C3MxuLzPi9mVihZXVgSi22OAYry6H/Qhb+Uk/Iof4jW8kAc6RFwDJNxqgK2Phoy8Sqjro
XbQ32z9gANR9DUIpL4cBxBBB/OJcCM7ciYXTZM1Ly9ZT0D7EaJPj93lFY9mnE2+kgcgB3qQBiI9k
pn72o7LQWg/zBb5ILMAtZKUih5J/ZWE3RFhkCaR2J+iqwt9+NhDR5PzQz2Nx0zu1i1K/boLf5Nd8
GB1LEPZvgVzuytyXmJOLq7tE2mrMDEGl6pBZvEmnV1ugiEIf1dpoWLc1p+5wGrOyaDb1EWYKZ2h8
t+48RtYNFU780RlE1PxSN1qSzg2pcE/u+SYl3T9iySTCB60vl/su//Ns2xQ7YkoUFtPJvvBEfN3y
HHJjJpyEnRUHKCksnDoTKJlwqSnMMNJMTj8jjVmy5hFigAVe6Id4eVmZnsudYze9HqGtPsDhopjW
tnrQ8BYLYpRRfcvHoxEeaFDNSuiidt9fNu8N04ofwSRtWFMGquzxNL8NaJeH2eVrul6Vbvysr85S
C9OUbm8GuDl1DEjBHTz/xmPoflpKTS+dRm6ECxlLZTte+U764yUZTx/s9wmepfKZgWudgkwI5Tl/
/nVCZxKrmB62TEZVewnCFxO+XmUmUfHe1Exq2a4/hW89qF1peq/wH/Qw0PnyuEcJ+Xw/3SeyU7vk
E/MP9zslyvxWVIK/SkVcIcFjW6x4hGQYMicSpsIsKLiQXts1O0kHF9RcepAKd5wBhXnZEZv+0KyV
bUlnT9jT+F8pQthoWheUIZqZUo0iqhRlwhRHrEXvOZhWnUcXtgIFIXPssZdyo3Ugj4ocuxl5Wz/O
oBiwq2YB5ba3eNSCarLppgTUARHAZPsDYbVk69ZHyBaHN875uyyT1lRgEA/c4f0sxNp6mtNxoi5L
j9o8pNMBcgJaWbA+KiZdB8JcxzEAobklfrqMC3YYxbrl7D412fbe1lzMG2LQX+Wt6TJFub5YifEB
o4fUcpUXwOvEOH2V58U9vuUEkEReekJ2XlOAjj9iHszbqN3HEIDE7WTmI0LSqj+Pjdzpmm0e+L0q
GSwWi115FfJWhziJaYsrPnD0ip/fU0EH1N8w5/yhRMOCDbrkCyQW0kWOqUBOs+DLlwR87eULzHVT
nVGTNsVzSRsZoNJIH5jsWnOuuUc0qrtKf9I7mDDWVw4RZtzbvrFVFNX56W/3VeyVLSBczBYPmfux
p0CN9GF0KnmBsJIOlKvULalzTNr2Hf+wPPW2mI39hSXNUiNHS7aTx3o986A0a38FKI39xiY8FIn+
q/KVKNxiXRMPqhHAMNFv8I5sSKAbObu3csfWXOzM2O7WS6NLVBVwO1jrBX3UMgXS+6IuLFuMD8MK
pWuIa9tzaYt5aJMmcRl9b5l554mtbIleWE9L3reHw5bVBFi/tz2g1Wm3hE+kdTufUp7VV5ywsfVo
jy4DnU6kbFurpYriL6G55YfQYyhPkm5Ifs8+6bsufNRj9ZvgIUT/I3C4BkORo/49ADw6F0nR1SPH
/PQ8jFHR7LaKio0M/F6d3Dw7vQvSsUEwsFurKICxmoNqHiTK1lXkI80h8g0dICPSlDykNCOE7Jnx
q3PUHqxL4pZ+STN91bDKqQ2ZPeiRI/cGaZpQWjTTGVCqkW2eTD/XkJ60qQUJCYZlylaGTZUHexfH
tBVwyXAXNP2YwKjoC/TC7rou3EMp46gd2kRwUSX8H99euy0xIpKzbleBc4OpXskQL3ZIp3aTjiuV
7dodUaT/ifwbSKzih9xeu8gcBhVmoEDgDefoyVGjVMPe4Hrh00383tLwxqGWE/eH0ok67U9expxS
epyg/G+WpjsvL0BRoiqCByu903EdvH5MdZrJFYp3F4stNgFEVs7UFeS1UkqVrMI9Ib66rIqtAig1
CjzW/UL5i7APgK4gWS0XTkWURZVuR40EKhl8SUBhpjYVzYtkxRgakcDiXHhaIoU0TFPjLwqn94Gl
ze//371RgstrEzkRhy20V58cVRa7XWx2usuSTCFuLrPeGkx3q84rn80U7IO0yCt+UGNca0UOs70x
o4L/ttLcW9vm4XyAun61ecHrVZ8eAwjnF0UhNSUXpL8LzbTUxV5s8mCC74lVzu9PiN35UgBQgTEk
MIslL8Px2OLFwXRx9q4wNKxG3oau0s20DQm2P1YRPVZkr+uN3XKXc9a8UdjJIYqUkN5IG9/ydR8y
KS1zvrtvaFOQuyvRnHw6Gb/eDqH5O/avZlKRcfE60RlaDaeomfK1ymyyvBh7zg923tV9yOXK8Rpk
EVTaVz4LqpfAFfUEniaXxdxUk7sD/5UR6+AlWOtORfTuKsooug4yIHW/YwsUPNIZd7o8vQjtd1CI
eK220c1IzL/nB3ShZaaipClz+1iuxZfaxWOP7OaCtppHYeqFAGERqpwr3RtsDIKskb/dwxWrtzbL
fMuNQBZh0B6P43sVZXDGWu4Ac9KPy9U1vX5RJzCN6oduzdVPHnBT6uwTrtKZUmKGBZQvn0CqNGxc
Zpzk4jyXVjXNaVlTWNqD4nMHEEDhH0fd4neVZymrD9jmVEzQEawrFzpXIn9Lt2NMfXBxZSq+bcyW
6h6s6hBV6cxSPvrrndbLB7jEPb1gBDO+9sav21G72vmidM8hf3MIo+wcE/UmHUpuLLPz4QykljX/
yYriAK22F1lGsH82hNYzny5tHPQdLdvMyioqPlynF8sTh19SrIedgitQyjbNn/dsQgLEI/erdPZH
ha4yxNHUJT29IKczr3GzxX8rQhUNctiLvJZCrUpTJ52a/+3B3jwuvcJ9mcJp68MzxcvQM70pWqzC
XP0b4iUs2PA7fuQmZK17fsdwIZZT60cnVJwvpFakjSfVEVUFvWRIPkrc/rAa+E71E57/ZCljR3l8
L5XO0z2dp9/MPcq9STmyYjgVDki0fO0mUel1l6OUbruXNXLYChK6frhGbBpN5O8YAii26mLxe87h
MRAeaGGJlUNcABlbGRBVDDRkBUchQCsXzQIml8qWucQm/6/8CZQRFrSEytDgnWvLaqpSLYPggGtN
lHbRC8smJozPP1peHdvHsWLJBqzyRNriqPfa5cRdd02tAm2JdyCuq+7x0y6qmlKdK8m6kM/Yhrd/
8ta5KYw5LB6zxcmwQcJLVknOmLbZ/iOmnjya3jfhZU8k72czd+dlulQxSlFzkr4e/SMc++8pv1av
ttV1pi1HgfatMg057KHJNmu9AL9vkY5qQqrbxAl1p3SwVbf1bWTPDrgSMMSB5QT7T5nuUyD6tN1A
fTLq7xe8jz32porS0cfK6j1kaDOONBd12D+nPAreL0v2bBdoWGIjLd7mUrM7H/WsuTE5Tx0YazBZ
oww6oTJzv/COC/yeyLe7UlVBLbEvuB2oQgrtR8GlHEK2WwprrqtSs/WfG33XHh90t+u0NLgRVKn9
spir7lz1+FA/vo/F3TC2zVp1F3o8bR5FEy4UT5++BW39uX2GkHJybdl3StafZCENXjuhv6uQznG4
s9NYKs04tntu4/c+voT+5YgHS6ee+XEuV6WWbFakVS9Tv0FxjxWPtHKu2PJc2miBAnOk7si6Fugp
0vTs7+XHjc65NfM8XPhmrOkG/d7705sOrQkAGgIRZXuDXC3nQL+cdE2tDs9/ykFuykpeJCTQlFb/
OM83bitJzaHoU14ajXJT32GywjBrc9OIOerLhRQzyeJgjkCT4GzY1jeymrMotR0MvNV3iv/Ti0CQ
bSUdRvEUf25VJSRcCSHFMdvP5RAaZDjRgePxW2VO+L6NLjR+gmQxjPVP5IGy2yJGKb0fUL5fK9kO
rmOT3DioYOrC2RmjEcl47x6SUqUajShL7Clyxt3h8yIs/lMhF/dvnkvLN02BM50SQLyJkBX9DxWT
uHMHM5zngH0FNNC1gVo86xHWhjJi011JlRQ1KarqwMCdis3uA0D67WCkeM+VIumUjgsOsy57m1To
77+M6UfEIkmO7Yn2l986XcA+sy7YCgVvNEztwCGRmqWOPsSnv87t96QRDO9yDI/VHbYt56NEZ39K
w1SEVK6fSJPHfgdks1x0oFlGwC8eOEnFwXJJyNs0hKw0c0WWdwOQjtoOjf3NVgmztqkVS1+bDizW
tNdBAVO6d3e4SUqEtvSDLROKbrmBYeMGA59KfqGFLJ3rBMnp2oL1jGyWxjDCLK7NVhpOfNeu5My/
s7jmHVnSRVhMbE8PJcelSf8udQuFeH1IPCRy439jUL+tSKv8rXxXh+X8Lo3G8hUki/sIfSdvIv2A
Y+Es2ulYuCoiNJfMUK5qi8s9O1euh2MaZVHcb7e4xa7LL7HEMNkX0XVQzCYbr55KMISi7lJvlcjf
E2IgJWZU5zDFGAHmxC2FsRv8SFajTzl5z3yylLEF/f1rIrf6p9tSTO2ZxB0Qh6uAaw4yufCjmz/S
l3IRA8t3abpxyq3VoBPg/n/huR5aoQdLDA6h52g9jjVwiTTi9H5nGMn1Z5/bkM/URUx8Dni89s0s
gkkz1Z3G9D1WiusYBxa7hOLKChOmCv6AV87M41Ar/o0hEfZ980wbgIpDotdXvzImtAa9+aRsq0IT
gr+sW3xKQqtVmtjoomv3zoSNcF0InPLPhzDZEEIAylP17PNSSmTpXIQY4D+6oJHBYWoYvltfOaaM
K0hGTNrFo+55YxJs/jkeZiV7BkXolJ9DShuRKqX93AqD49znb9zRxKgK1Ycfw/meZA9s5CoFfiEE
M99yt6BzxAvPnl2TY9PDgmhnk+iQ3u9ojrKwVh5cwUpdPLIB8AQ2RvpdqYSrKPmjLzPkhHks/8P8
i/7lq9chEwI8PRVaAOCkrcXttoX73TegEHOUjVrcElhvdimdygOppd5P6IWGaYM9xuQBBIQAFqrY
TB4w1g8hnaKC4o+rkqP5EEkHbJxUFgHAoIF4OpxwUbADYsCXPq8CuGGqGHzi19TaPWJvC333HU0i
eJbVkPNbPjoNy9G1gdWRgmD11A98F5bF6IDZqjqdZPiY8rSLSgkI5uWjsyYzr+IaJJTiW8yKov2R
obsOoaiaK9WVrCI6fzjeipqla03tmJefVrBM9mJJ1nPfb0uIJnWDY4tmd9iu7xqSURXn9vG8dh48
/4tzclHx6sh1YE3e0Y+h6YgQRCit2dD/8VPZSL3GA6BMyC++YMuRkEr6MmuPhFC2uDxLtUPjueuX
MWC1eeynrkVB/naSQAXY7ucm/Jn9m5hxXqKBKjeTl5w6mG27qAn2duQi0UN0Bzs2E990VGLz5MWQ
xbJZTk3V2mdW5L6a8GMKla/+SWGjWrqPDiVXIqNog4n7NawE5LUBjuqjsRj4uuncas89jVvwTlct
+D/yMliZVAfL6D05fUbD5Pi/VCtvnoYPGwyih+TijJ6bMEkfRmyJKyEbtlM1rusGUnGizMMY+tW2
/JUjtLge1yl5jsbT+zZd6RFOC7AyqFvtzev4bhONz48TluJzKyfWdOk23AmCdxSYmVO4auRvlCKf
BFyjgjPmEE3oaXq1kd1p/aFWgdauVFxl84ramuPIgRAILqloU2QiyJTR1+HTlcq8T8tp7m2cRPMA
+zRzcccMWJilbKPBr2U6wqoC8kXm5ztSvLuindCx/aqMmxlnFnCsKqA+DwWLQQG79R2G8pXuPR3T
ZjiQrHOuiQ63jCunuoA4Nuq6BRcP0lQ5nqHHEhKoUhHLI4omHRPGva12LuNglRfbrsWCYGn4VhMJ
vesTHwUZi6bHgIHQJDBAP4G4JDGVD8uaQZeKNEHS0UDYThHW1v+tMgie4hVhtelrsowpYllSqYfP
MbPTUwdX/xrE6Z8PNT42aClbJNv5tLlFIYt1g97e82Og3P8vyU+62Xss5o+b4AQVTI3c6Hw4JcpC
1IjraPTRAlXoFvBTtJEglNe/MK2xln6fFs+iRRcOueVIDV21WHXdQ5oDpEZ2dokpg/7psyss8TPi
LNwkVxXr5W1lNXyas5OGt+MAK7hHqxTVuXK0W+g82Xom91LjTn+XKXTKmwNmqQtxeIS9bjVPzu3J
ImSRXxmbH+DkCai0PekjJGpVqpRTi82GytUkOf/KqPnjBsKIXkCxzxA7AhsHk7qxaaWgznfK3tr6
raSa6wO+KYIN/NalSIyeVUcdrihIGJfE9mMrMnieWLIc70PbMyaxc91lv2SXmr2lQYUxKXcA6o49
6BC8I4KzIIQ0JIx96ZUyLUk6GPUzj0zX4ClbKlrtp2d3aXyWjo2l0jfTKfy/aMMJv4Z6TfrGfEGL
cCFZuH+X27QWmEPZdv8sQgVbVS5fzHgaegFWlIGv9BLpxi1bRhLsoI5YG9E0YGEaGJ7hbV42Nu+l
0GvJrYqXICGWnAMOFZY/vk4xhc4XaXgPm6OCEGC803LC6/pyNl2libMslK8rrqBpldMpdmfHTWtI
y8Xh5XXVfxkk4e90k5DMk6so22cl/ykn85XutV5L/er1aypz9pvCyyS+JgkpiaI3XF/7FTLfKLt2
LI/XT9TSMZ9Gbez63hgb0K1HA70EzwlKnCg84MvZc4zOP0r13ey2uLLl9bJG4OoQQuh0F+Jr7Dcb
ultH/9a7tBa9om0syfGk7a0pwQe1M9JuQUAOAhhMEeMHmFicIIngJu/TeG7gMkqGJhfp0pxJr7kx
KLi1qiqfQf26eXLB3FSne5+kregMzzkRsnSEY4a9w85GYIe4YoIYQZRHD5KRNR1iJL72EOS/MJcQ
E6igdx4B2M1y6BQ2GnydWZjZMVMcRCrDOZHvnakcBP2M8O4GYkZTun29L2Xag9P7NMmT66LVivUR
B+LQ8nCtS/jYnzx8QYBuccdCVfervV4MKMXvdVTkM6EJRR/yjJEx4d5ICtXXAjpaLhb5TXu8TRvJ
7e3kMl2jxwf8yGAM4Iz9U++u72P26rVdcLkKvA+9Md8pGBmdTn9N5Q1xvvu5avVQO/Nv1NjzBXGY
IUulLEaU5qDxAJpKFvKiMoHhBhEetP2sFOyWMwxgXwl2p1ssWc/ahRcJYyB9GYlZR9WPElKeGvC1
fZIEqhrYgPCwxbwJbi0pcCpVtmJd0oM6bS5zGgQMmuJ/X8ocRYDZs+oLc/GTjwmeH6J1ji8Ew4Z3
Dz9J7pHUCSX7YF8RNo7czhJFCEEyRdLqOHq62cxNegz2i+TEJpxnF6jzaZHi0twkgn2N8isZUJEB
+0rj5QIr68rCArk4NEWh5pq2mOaLKVUR0+B3/gtwMnCG+ZtOjL7oYYY+U+S0n/M73kMonJfBr0Wk
XaZRM9cQKFwMRpo5miEU0wiNslTQ8IO+hJsMzUnFvU7pZj2rUXcUkpzDCTSN6Vd41leSxyvdkx0M
8GejBr8/9tNn2IwD402fXSK1G43q6TxRivlfss84xo6L+n1Zp4EOtE+xnWUB/DmYvnZAuKAV9MYd
PITcK3T/Z6SYGsMq5ey5mQTV6djZdUfjVVHz9MwmpN9Ouzh3AaNC4Br6oFplUmhxARmKLo0k4bKK
CmnO3kdX8wCdRZrWjDxrCeaxXRuTSG7mi2AqCqVbgasxC8uR875mUdlAUPBie6k7RVvbFWrsEu/n
LdKXLxaa3f2KuebwMDiq2RbOMwjDgeNKdi/ooD+220k5R6SH9A1HnlNo4pIvYZ2F0nxBNsP1HjNl
r871twYYlJy2R4PTu2w4ae7/imK0szBmTf1PaeTiyQyclYAXAB90k810WAkh8E4Wg2AZAbi2ninC
ibfi6niYQPlRTUSB3xKQg1EkcsNqxQFSqNlmsrdL5QzfuVwCinmi8Iu374ho36PDZa+8hn6DAufW
UccNUmnk174O3I5Gcf5jUw0qwy4QukZkcI1zJYTIntciL+47ZSewI44iZVynokAYqb24zsJYwgdm
hioUJWn17M/kQQdUisipqUCCDMxQs8CDSzIWbkERUOj5U/f6/IIGyt/Y5SxbZ1Tfo/v9oTkiXGiQ
rvEzt+sl6IaCGHf2uCBhY180K+aRwy6vBJRctfUXeko9YhDWtDJ0PESPS4VcCv0onHWZUjrSWGCI
qMIDliCG1Q45u5ypJxUBzU8TkCkul0k1Eby1/TDtjgD/zJfTi6GZMfqHaCYzRB8ZzvI1pi9e98Da
RQiR2gwfSVf4zrlwG9tgmj2QtCfT1go47/RqFkDu3oKD/ocOzZyTaZFtlVCKpWSr4UM9ghZ8etNk
eoQRy8koFbyn5vu8Z3fcUNChoCK0wmLqLle8QCtjQJn6L6DaZxxIo3fEpJTYOAIR7nAfcp2hOyj0
oGY0qZde73yyXq4yyYCpFSyBVZjwlg8EobzcE+Wk9HxInQAMvDSPipiX6j7cyJbkZnhu2keoe96a
ALMcUgMLICI2LxVQam/8DQ6SYdaVmmQWge8Gwjl1rhLLoobkUDSkZl6S1DiVizoSiz/Wf9G0pEJZ
5w5ouD0Jfbj+Z2gfBePtIIukrRgEWCtjKQ2p7qnlk6Zwjn+8xkGesog301ngPQLjYFBllE0g/gmi
JCo8KwMAacOc0bjl39Jctyb6PPNdFMUm73Z13wRmOOYyK5IHJY5hk562zUu69sPWDcJUpvxmx4hi
+R/40wJ/8Pn/e7Ji9nxK+/f8EyfrQcCyrSxYHl7FlkYXi3KGFkN1dxYSBuqtvS5I2gwQDpABThhV
NakFORbncUrpz1+kO93Fr9aPwrlQvQZdvkkZH02a7Equ4O0FAPruJ04sewEztD5X2JbhBSyB6VPM
nRdx45boRMgtEsADpZkQzQniJ4GevTlZJNJdOp42xm8vTNI2wgMt144ruhrXJm6uqhxzRRcsL/na
zGRmKoktAyCYsQSCpUj4gNv6uilU1DuA8g9ztmmAh4zBCSBFAueO3ijHyFec5jpRLvp9TThk65Ot
N0vdUn+0Sz6ItrzydqY70fAQ1e4JKgBoN0g6zCL/oW4XKZ1zH9DffFulxIPx/XUINaFkKuqG0ECo
yBLl0CBVP8tjUMhnOr4Qz6VT8KtnlhG4A02uFv8xHmaauBAO/FBRO1aJeYUxND2bwNtmDDeLRtPG
psk+iTyDRH0ijBJ+KW7uAJPgxedXLiFKd/dM/W1PGym9qgxQMdGOpP4mnHGE9NSAMhgaLulkpxjZ
gZJRxbhRKJVA55IIfKlK7r7zRjoUL57GHHNECat1REDs6LJukA51b3pc9eXFfQ0/OBl7vhEh0tvR
+O/pT00Xhqnq/adQY9MvzVca91/NfxmjUdqYIWYOdAbH+ourmVvVmIfRFGEeFC5ixNDSyFBxy2hY
BaQsn6Fu5Etq2UbvWKTIh8DfwMNA3MeVqResiz9pM8cc2CYPiWFndaFlTW+6ewh04eLLvi+5k6mP
FCUN1iajgMECHsT03ObWROoJVDmUT2dVoIYRLboqdDHYqHrNSXtxqB/crsRjdc4r008oLFBr15ly
LaPyZg3S6+yK9LTO6tvLvud9nMcNRLzQKMkDx8ChQ+ZRkkL4HMwC0KLRVDqYbLdXuHugHddoPSkB
cKmNHquxh3tXMaamjQgp50c1smgzy9okhzMfRZhv7IucgoGyKk4k5cTFde6aZ4QH2XWvJT27jAax
1EWwl8oplXAhOr9n5trDbUWfxVUN0lldawTgv2MBUXBcY/A4PRR42+u7Iz+sB37+rb0dVB+iIJYm
xQrn9jD+dnv/D/CIpp6aUETxaHlujLy7dR5iE9Cmw97ktErNDdOxIUl3aCT40Rj60ogMpLbmKZjq
TqAH2wvCJaOYckYH+L3Nm5SbkpFZOvaOnqd8V7P11OHl9u6wx5lk/3IwdOOmZRm0Sfwc4A5vaUfQ
wuStScCjS1gr3LmybpVhXAjUvHwFXvKQhisYwmphKdEK1TVIMb6GY8EVpcwrn3+puVCSvspv2QNN
X+2ZiwSDVwpFHQxt3GKFdYWa4ib1AgXqJU14tKn9EtnJs0JXsnmie4u79GddXyuoBKr94DM7vkjS
o+cmJ5HYQN724zWm3TxzKq6X7wov9tTE8VQmxjOJ+kI91kvoOoBvKRl4yQ5tgcdfAz6+Hqx046Am
Fu+qSyCedg62PhBhVT5HfSP8kwNJIvFW5v9k+BjhSDgbC6M5kDfi12ekotZX//0Yumizmc3tcBMQ
ErSLZc50ppQJYBZ+StJKznWrH+n0giBko/9bGLpXRk8N5ICjEjTtuitT0+HabFyVFDb/U37DLQp8
O9ffHBamwlB1VKN8vgCF+3I0K+nWJ/4fi+DJneHT0iTNvFCFucp2eUpmawBK/+ma88pUmh0itrQe
L8dEsTZoUQ+kNKj/Do8Kjisj81OjspriE0ptHLs64fVPJlkuCfJR7ww/oGA2iSc91MM0l7rurErC
HzUHgLTwJGG96yWrrh+PBHhjU6rj3/eKdNx0PAJvZgswIoaASrHetarr+OQKXsqFkYFXvZqwfJ72
wrER1O+9IaVRdm3qn2NdQQ+8ZlTbVbhH7J6PZZzMQmGFICtATA8V5vsF25NJL57L9BnIpuHSH2g7
a+PF1RAveeJt4oLW+rtxLMlHp6GeCTYuZM6pJlyXTpMsuGaVRjbguYL/meeo77SIPY5N2/zP5wNu
lsXB/kHc4ng48gL+bOeyw3b/HAzJAqulDfawxQXYXcqGN7pOjt/z7rmk/4p8G5y16F/tGby/iP2S
hqYDVhk/otnKblsM1UUVdkn/oSKH3AJfH/InQzlaZSyrOjnBmi9oGE7UP0gcvDHJ/Tq4IDx6iVf6
rzkVOhhgteSdqhM85OQA26b7Qe6ImGYiQ3SepkiAQGyAiMoxQiVLIyhLMXnP2yx6PgG43jKEDUaW
k66B5FkKWrdX7Q3AE8IzbB8hmLkUpOO7iM4OGMYwRlbLeZ5ALG7Kf83vhO+mQzB//sDIOf5cSG2t
jzdOkLH9IKtAuuxAShzUsbA7Ic2+qdZyIubJ/wnEFNz6gO4Sleb9SmH6e5yZ9XUSIJDbHR4vjim0
ZPzclcbTgD6lcJ1uKQq9Rzl15XKHTj0xTtd/S927RTPaaLKd/uT1D5PRfDcxxy3odwxsgtleJRrm
IZFqJy/xuMu9CJoQTHe8OHwXWGG+NSaJYZ/N1UdEMqXu6WzWTG8xGoB499VPGEktdqfvAxAHLzKN
qQ6pDLnZX3cKo+JgrFJK9dBYavxpIX5hOF7wpglSYXh20z2p896mOVcGXerkyx6zU3w4Ik6Xadcj
4KrkYlIxZYgD1Hkdt278uBlje32q7QytyOfX5BH17XNES5YS9qSducX1//kt5bHIi8hjWVyRSCsr
4qWE7Wv13w+7xUyHZIkFYcsOk15DHtCf8G6BHsCHmPpPaEOQP0eX5losViINxkOpIItdi00HdJ3l
I2cwFUU2Y17LiUyOJX3xL4Z2xEktCsHTpr2Np6ecoXqyXmnMFdT5jz9hK6rLRG7xnwQDmbuFkQ2D
ohZKJ4hYfSTqcX/5TvtdgyXsjZ5lfS1h+7MIApN+vZi27OG8pfRpk8As6W0ADjY6rYePRadyVBdE
Ks+xShZ0grISRL+hcKUgrMNeEudYSsKMd5v/Mjito6SBLoxQswwhth+Vj3wRst0oBPmlO80dq8B+
BI2yGqWADFLR5nxlM7mOKnvMmiWlhDrAWXWDmDtzSm+A8F0xD/tH3Mqu1jV7sfd865ACULg3ii4o
TaF+QYteL0I7cN1CD8sIlHNgE8iuuREVL7tmzvOcx/4Rj2BUlhLc6WAqDQq9c6DD49mvDsWabaD/
/poKW8fer+C87zJoTXHcf7nMlrdEz7ZlGRmuLAvy3VLApxVAvpM7/3QepYCRSZcNxv7JITn0X2zu
3XdeNklMSwnnimkHPVCkEdC7r9I5ZhKPxy0+b/KERNut6WQ9BPMP9vJdvRjS7zzXiFx9PeKZvM/r
EniFUR6BHYRMsOl7rcx3H9+PiHDwkWRmy2v48iCyJM0mrI23X6He7pMTs3+bmemjEJSX0iLlud8U
T2WrPIO14b5YlVCR2kiDBzi7+9suR0zSGLQ+WmcJPOcDRbmYRZFvF4/CZ+OOTYHGNNkRHhjJoD8V
VfApG0OtEiCr3bA35NJ9k7zpC6P/OZa1Neq5/SGAj53gu/T0Fnk0wVzULyyBn6vyJE2mlHaGLGLn
kCJuETvmhp+/6YgUnyeSqc7ojj/7JjK/C90fw3zsFmbrCzU6WM6KFrhRNNdkSENLssrN2r4cR52I
6arq775zc+RAHM5JBAM7/cJ98mCFsYC5tYtC+kLEnMD4VgxRo0ntb1RJe89icM/2EaKCWdNz+4lh
1IbIJyQ4sEIGmuSSgipNoIdvd7dN+Ew4jd3nARW4A45Li00GOagKgx8F0FUPP79zwT+SrkJPdMg8
PyfHS2irvdjDLwsuomNcM5/JYdqxLVnlDmDJZZpNvx4I8EJqbHOzp2h3g6/bCQHIaWt09qP29gy9
Qb/Kq/Pj6a0U/d6TuPAxDDGgph9RLIbgFK71jhH0IxSyE/TehOYl/wi3LaO2Qx5PXLY0x9ZFnsdd
6L88lLe4E4D5NB+X8jp5RQiLLVsq66SV6pbJYZQo4ICZo3J2b8qIf0782E4ABsI0Np0GVQ5fHtRq
HUC3Dy8+hKsZYZISy1Rud66EGMFFIKB5m/q3zd5Mb/4EU43D0iQGZNrUq9dzUk4pdx0ezbAsvBlD
i3fWMAoLqoVeHzC7DG3J1xqaRqoxpEizg1HrfX6Zg2bkaS1mHp+smNNmKkjy7zCinp5HtTmofVyO
SScEhwBHQEYlRqDEB3jT6rMZwyEGD1w0vMhBbK6ArvGq6XvBgzuQX5eBspXtg+sbaQhg6/Yf4M67
h6P8lKbvMAzHnoZPKGtapmyeHD9hw5We9gXT6GTpPa0hpBYu9RN8UKRJMbqnDgTPkEtkGcwMJdbP
R+id2+7XeYQ+wSnPxgHL1PAHZypSTF8Skyt7Ncao5e3hsg0eZTgkXrieWGBkG22bhDCNGDSS5xVV
y1mlvAjtc2Q4sVIMTsOYHP8XTB5JzTS82M4DkbaTDWJ01dD+jG1Cp+F3TnqjYU35eWKXz0aMQJzn
EL8DVucAJKXsgubb/amltTVkoZ4uB0eJFmtTDNPHt8r2nx5J9re0TBkylK09t5ss5Wc3J0jI0Pet
zeb34k4W/x5wVOMA+8OEZSuYSD2bKrkSaAN4PAHymIoLDtdDjug+8KObwQmyv/iCiJgjtrmB58I+
m0BKBKFMH5Kvbsf214HiYWo/OGjWE1gTtb+1zwW6xO/j1p719RIRmY3r2saXMZz+XqGfgeKHufDc
9tju3Hdd2maX7RzO5flNTnba8O3zPpv1IB1DqbFmFvy+KTkYqNJCKdjTqWAwU5f6sPnLTvEuHFUn
cHoLjIXZbZv/nRNALRRF1CPlCvthw+WlfZgTOoZoAIfGy/iJl4uq1i24XLpIqNx10wX5dhAgUMyb
tEkhnrWBLt7W0sOULVzl2URmNWK9YAPvpoDTt5dP1Zsmkhv42iijAGwLkujSWsrHsrhdYrXx47u7
XlkTYTXgut1IWxfOKDGlaABI1pFCejCI9w1AvBWNILHI3pDU/sTLsXKuNoFBpYymtm7s/CBmXzdo
lwRCmiBZK2lxUk2yqVlPJl/A+G8oJECsjYUnV+o5/aei+FpRKOmIoxsJV+yVol95JeEU0f2myayq
9sjpZkI3nL0axrzktvZhazJ4DCQintAyGWGQFNaa/yAOXyUB04H3H2pWnfCem2ioMU0fa3d5MT9A
fge0rsLAnJkyvxPucNPJ+v2ukf9+r05OzQPVC+/2reIe8pugsYPQ1Gax2zkyVa6MSExI4YCBN0du
XedRxT7hyBr3NjlvpPttO0dTgNjZCILo3p8S5FMFwdJjnwWescdJRh44m2pb25DueJjonVZXi0qS
77wXek8yqErNt2zlpSOk6FqEV/FdPWc5OI0veqU5FOkhF3eToT8D1NrPs9NWP6D536qhfHQahZZ7
nJVjjBMemlO+U5WPwQv7wau5RILN7xyWCcKWnyxLbMyWBc0oYvbHxeN/oVjXtV08u6oYgLirgDRV
Rw/CPMXAf6BYVIxvxc7mfgyGUVub5XEFYdkkAaFvJxa2AlMsGLo117drq/1VCitOrd2jeBOMrV+L
FOum/ddK1TylXFufMgoTIwFB8AMyOo05psbyBUswHoJqjwURRcOlMAjKlwadnkF8QINBxs/z7a6v
NfYHm7hG8/ZSO2mB03qtQN/4tRIoUGH2qmmdWTq8wNpCxIXXhNg0StrdRrNPasBW1Gx8r9gR9vcB
MGoDrO+37yRaomTLo46HPbiP3TiW+5i/JhqiJLWksxJJ7FiJOxelQdUleX7/s7QYGsbwKVyUKDHZ
Fb+M30XrPrXa6Goji1VPFJIpw+lA8ahhJkzkW5M4PGNcNYWgA9qTUAlhUJf/tnYDSiFtNVfIAYp0
achThNAzpGG4+gyOUa9/DnLtb2qyZ/kOQFqi8q/tGQ9eRja6dgU7ovguhKKxwQoMJGk3GRBhfDY0
bcPMBr5763hRHrV2Sw1Sy892cRd0MmjphssvQkUCe1qBLK/7IFLUiEDVoVO74yCQMHDHlAwBSkWL
xeeVhwhL9xrwj+jheu1fkxvJa5Nuxn8nAzAFQUKkV4IpmP6cTaNK2ThgtDmjG0EivXuJRjT4/yJs
Ykke3PXACW5MEx1ZgBscfXlMGScPxY9nLAeOGxXxrY+mDnFJGKsyRWDimaSQEtst5jVenN0UNw0K
/rjcMyn4z3dDSKLERjczj0dErdhstkKOVa0pkgT5Gqf1LwiPXqO8B+wkPodKm6oMpehCSMMggcEF
r9jnUckFHsoSKhVELJUGGW67fPHkZUcve/V78asjpEw5gQzQKvtRekq+xP+6Gecml3HNR++Z/FFL
BtNjvGKwM9KNBINrveNaCDBzGxAOFIZ7UmThsNt2qS+qZEJLdWEeQDrefOR6TkLxThHM9sK0IBj5
ps1oj2e3kSJKozllPXsXNLoBF1XADCe2cFLuu+R/0uOKJQAugwJLwcnkfPR+6rutlxvW3IxdLjQX
/+Yu6XrV/eLfnojxstDxCRxiy5OPNhGvlEHhoZM6avKHUSFCTppvD7HwAKe9cuQceFdYf4OStXPe
MPzaTsxKnCScuvKbxI3qkfRe3u06J+3GqMguQ5hQxm+Q8neooYnAAtfP6HTKXu70EhM7o5SQeTk4
eT++Tc2YFCalV+0NRMiUOcq3kNcwvneRxA7rgP1igGe5EM994VFhWLSMEkrklz062p/qjgC9KDd5
NQ2neKpGKrhzKpC4iUK1Zg6p+GpBbNqHwvzMerEsK17TrRH3xamgbt4GYjyn9g/E4r5Njk9UXGZv
set6hHSeOrxy9zkBgInQQcqwP6PsWXrACs2VN3R8MdX+EFsD/1O2u4l8FxgjZ1t7YUYpctB5tWsz
tnN1EN9LE/9ugHlliTfAwnzhS3d25DHJe0SYkzEU8f/LHFZAfTmwoo/VO8TT/L7iPTk+4DHcEG7U
nhr+NFmAduN/XYwS1SadFLAKPWXS8xLtOlIxDKGzAaa8nPqqhXEf/aziRYG0z56WGNjBElmkemJU
TO8Ysn1HsT8Z0hII4wxbf3UzmrJTIy31YFudvpYe+UcybGmdpStB8yNwZVUSnMflgl8qYHcwtpFw
LKDrVfzWUjVdqgLIGrLlFMk9e45+VJSsnq2jQJ8vXjouR/IeGdYie2PShNmrPm/8bUGlA8cK8UmR
ILoUKaRP6QrBVTarsWd/dIFHEqRjpV6NCl4YheyCp+83/torCCwmE4/ZaIBO0mtj5JHWdaKi99NE
Q/7z7Els8/l/6MdXWpcuzdjNubL1+FgKOFeSVYALcVf8mjeKi1Cf8vhhUEeLFSSQvZQXk4B4XEEU
GJe4GUyr9Ap9h22oQaE6k3kAR6rO0aWgyEbmxTl4ZipKtbOdqUd61V+7ZzYwGZMCv7RAs45lDWVM
7z/pUnV9zjEClxhmw7pdjugjH2uDjP1s0Zc0ITrnfr632S1EhIs9tvYFkFm9BAoZIjHxL4ofl1oc
snfiV46z7jsU/bgbYgGnxoK5RfBPc3JlK9PQkwCZnhGrCMdBkrBZb3prMMsXVQf1lgZFTMXy1Nwl
MB3CLuKBpG1Hxy8eEbCTPvePejd3Bd4e/MBNWfzetjrGdGU7c6X116LKW4GzIaDZ3kJF58RiUPnl
nxrqLstQ1D3HhMQ15o1l5fp3quuY8e6Qf72kbz0SdhI57T/xYoCxGWlcaIlEIZjs7Fir6r8e9pqI
OFSni+jQIK6sPqgBQqan06DgwcY/2Zzum1vgpe4OvAC62pdyWMzMkfAa7eJfOeeQ/8kWU8Ayw/qD
Dlpu72bWYi2qB4VHEbW6jk9MZ9wTFMfK9+3cHKAOwBu0XM74bKvm9/AK2EnPpLaS/y9Se8AX7Kxq
UIvcVyKzmsB9YAjbZqxwaMBlsY4X8kzzdE3WTyqgbUKXmoDImdCwhzlVDyfmrOZoYyr6JJKG06oB
tI0WGCJSqcLwxjsfD2X5eDu9HOkSWypUJ/dtgLtd6fsqHzG7Y73xPXEKtEXIgkyHUAbK/TeeMKNa
ZUaFzWYN58DAKggVjlmVqxotNTux9h5eitFDGZ+dXV9E3i17KAKpkeXqKMxvhOw3kyTUXlK+lBQq
ugtJ6BCH+ztxBwmKMn9UTPZgrfw/QZdmZKjcrJhhImOuWgTdK400N1l7ar++8lZIBO3eXC1XoQBh
6mbMf+X26nhHjPVrTwIkzNBAA/Q/oq5iUcKjpvA8DabQIdMhA7lgU8cz8JcfMp2Y9h1wmWWcjrhA
Gq8JztkyoBHHBkqePCn1EOtSDaXImj1xVTnlcTYxv0OAs/6UCis3SypBm2UD8xbFZoYerzp049Y9
kncNsAed0q0aA/yeaNHPcVs53A1fN2V0QZ1Ao7INHDOMfyKs30ptnek6wMs2SmdsltnLhoHNlZeu
gNm76KXUPICyL7FUrO7pjVsKV6ombu2+PMg429b+d5gxLNGNQgyYV3aSll0RC+QW/NzcupnQsT4P
d4cWjj3gSK/X/Ao1cWH8+N3eGFfWkuzLH2EHsiQCmbVExQJpdzDbhSi9aGl+PcEZfOQ+HByx3i8V
ZlMDk8yC9GKcrxooQ7r2j7iYBuESQGOV240Q752LpW9KPlge12R4YiAOsNWrhxv9MQ/5vPPXg5XP
7JWkJP+dbWTkRFbfrwsHS3R24gfOW7Uq8gA5DVgQX/FERGaH+UDtntgee/UZRFvIVr3i6k0QN5F1
zU8OKcn0HCAfcu2b8/cAx07aGV1KT6M+kYfnGFpOoCzGS2bThaC3hSC5vRIiG8G7KjWqc6pqgzM6
oHX/CY2wCG64znrdy10j/5Qx+ikKa8O04kzr1Iey8u+H2u9tReNjFJMmvbCOvAwpECDM+8eiVq8L
8Dl9Clc+d1L2VMmQrjUpex+WLMpNDZ4LC8N1JQMDcKnu7WMMRGjvyeCoYEXZl0pK/6YaJyCxpG71
7Xgjtea4Zq5zNvKx8iCaoX4LPnZ1ze/j4QMJubhcWYI8UmItE7S7XOKoChQTUyF1yLkhpgkrlm6B
oOlLv139A3eTk4lK2JYFZdRB8T1HS1x4q4gSLa/X6yOmU1uZkdyAtHZbPccWlauCQWmvDutWkl4e
TiOoTJkpmb4rSW9IK0TibsGo1ei2T7LH2LJq/cXbtcUidB0+8/YCwqyqqRx3SsfFoRrTV5j3hf7+
P9qc/o2/D8k8l06bVVL4I3p1PFTanXDcH5TfIU1meQM/eJgKViAIki5HHkvObF4CtBQehyIl6Jb+
3Gal6hvwAgm2Y6uh+h+J+HhErTKlRKMXaVHnaH8QVed9tUdUah5uIyTEJRQPG8uFjmzdGc1yblKE
J7sG+od+74ol8TaMrjQq5TrA6nUpn4hP95061Agzb78lIKbDzmIljQXvYURkxnNK3jNW2zcSdKgH
b0ST/ZHC0Ymh6dopEKnXYeK9ullP3y9bHzYXp6UwffccboA+Tf/LzJgkGZ0kX52kCnnWyiGUcLse
zyVX5ZECkGv9/QX2GtwiMLXFyKuDtL9aVcKXVjZTPN1KsGzpuRol/peAvjlPleQ0Natbx8MHhbQO
uyP1mjPGLGKAoUaJySycSZI2VRfQ/7YEXfTBs3QCPiy+g4oJzHX89snNRYfqwjcWb/oMYjCbAg/9
+OvxsE5NUMhh7oqlS0IpUsqj44wuGfy6OBVPptE8x98UqI67j4PYEV5yTuiX+ANKdE2QbWYEzp3K
9CjjKItfK2DP/bcijMBdB4asp1wesrFQj+CYVozcoFzuf4wInZwyG4TXEEcvqekK2H9JZM9S0c/S
OGlW6AlXo9oV+TdCv/Ylm3ClAEcTN+XNFPUZ8b0h0buSGBpwun55evIEzXzYUia7nO6Axk62V50I
Uq5KcHANWIjl7y7xyV/vT7ICvB0cleyRhnLu+I30gA9rTkjUyBe4UJRJSpSpSGD9vnEialHcYJKo
YQxGIAIZSz+WvkmzAWUSv6X1tFK61XEl4/lI6+28F4EVgLFDMtsIZ4/RbP41eGurk1n5b67mXjSE
lR9hp1q0l3P34AXxeylF+w/wZ3+hhLZX56ZFLQdlzshK1A4GyAttiZyKakO7LdloeVwF6JTmdgq8
aEGw8UyDlRHUB6iH0mcqKq7eup2qs62juFbHk1MkTv2DO9kiTh9C7UGAZg5gAll/6Q/TC+1TLSdr
sLAU1Mk2qAFDy7eLGgUOqUD2tagluIPM1Ti7M0r19q/XcDClh5ZvxhKAyQurp4w5aecb54/uhDum
KXA2hT2bW+n+wc4g5Wwi5FGLrzyly34Y+e186RlzRir805lh6SVBgDPZOr45tZNC9ytI11Yi12mC
lsP9fsJ8cQWsXbugHMp+wPBwiJWTv9S8z4fyKOSExBEzkIgE2erfCnMnapHj2JS/jPU+waCPbZ+6
DQE3SbZwS3fYjdMVpqJQGnEl4gRCcvRkMYM71ObGVE2VJB2FBw9i/nhr/IXHeMO8UTM1CB5/xr/N
12bSR9XfvITw/ajo36YcZS8CLtvsTwN9C2ZPCk2bq2cyz5ArO1U8uyigKvfr0Ow8jIxm9ndAt0fc
2VllvWmb5oUzBNZPlDMvq0H3WGKEowuDYD2AveWPzJ9TmEgtx30zniw+SCgJcLKcVF6525rT3JNL
WvFGJJv9HyHZd4mNfZdIDgcCMcIdBgJwYTee38Zhv+Y/qfkOvZzAsQyWlJFrNAKTdnzUBIoktlTD
+jiqBM3zu4NGaXk2ndHmNRCoOLWdsqWQdnunROBlVgIyERW5qx7nl48PWiExDzvUOJwcrxmF4sST
04H+RGO0icPBDPIINT5rtR7VFzdh/NXBfGKLr5+TMKx76NemgRcbhw+pedJ//q7eRDm06i4GNLSh
cmrJqONXb7GbRCPNbUBDEId7l1H4XK3QfsWas8j+3YkqWhbZwB6W6Hq7z7xB2guv/GElYhYHCK4t
hX6DolRbWP/2gtGnNtpNXvA4x61MxIOHd6nTd4XiHY3oszrItPDJuwZ/B2ya/wnRrNAFFYu0lB0n
jSy/Wd9AopMTLWu26/6BO1broX+XYfTibQpWfURfGk1B92oD+VoYv3bXUDERCQ+viHbB2rKVgiHX
fxRztSogq2pzhzwUdSbKP2IJAPVGY8VoPlx7ziceks49SwWnV8u9/BNxHXC2IT0ce69AjjMdunF6
xvcfRP0575wSLZgOBLhXCxDcCvzVUXtIrsk8SbPxOcfpIOULOkDlCS65aofh7CfO3TSZYrbywsY1
n7NLOuwCTBdouzx9cl2wxntK5H96stm1PxOp8xQJNgZcgXXrzOPNjWyvfMoO194j/JP0z8pduGiY
69UFNeEvTW8U39yv+xT547augckIuGpZ/F0xm6g/468o58r5RRFZFPL08SyLQzV2I18W+aG8rjF1
THvfAFCi3FyiSGtjv90wyKgLBALYBIT52IGj3OCLZLYX0FrSJ930yIhEcuFhGTf1AaNNcQg09TGV
YWr22LKbsarK5/pe+5QC2A637PbKbCCrOAcNQZATVnh/uHuiybQF3Ud7hqngxf6xKC+CvphressQ
jG2TDA8xa+3+tZERqVbTV1/F53yuZ8fYTARLLKqVxRQGUwfrDRcMQGqfbOmyFw7/VsQ6Tv/wfZA/
iJVnLgYEhK0jk1tIJf0+UaKF/RZrjVpyHQBVx2aYO7y74lqLylktsxFsUb0dSJkWsxCSLzDlS1Zb
vJVxKLt2WPRuojY6mTzCWzjzTZY8BaIQlMJ1rUP8lu8pvbMer9/1cQpxl39xGB4fIrWVIlejCmQ7
xyjGIyvCTbb23GBv5I3sqHXZRCixRzmUWMe2++ULNAM0576bd8w+IVeQLYa1m1liaxs8trTzUUaj
CEJVsnfCTkj2/2hh1WmM/kEAHxu6A6s4aZ4htEpVJ7C/6P3yqpcyxMJ/6B0MD5vb6nhx8lZrwdRe
7Bh4GdJAmQiKvNn4XeJV+sJXfwwuo77wvTJZbP6idq2hgdypOeTGm4EsTgzrYG34m/l96dglcLyN
4tr6YXPLF/uf0v2CH8rCeJ0kM7ji+iaHOGV0lIxXvnUFQf++WU4BBiV112w6KQm0axXg1cgiaxsJ
TTscBnKBYr49hr5WZsEmB3GKKdHnIkjZ3zaq/vXhn63RGBrHY0Npv37UtNbsSrtb0upSEMJQJNIB
ZGmtKbI2Eeb5zEjp3ROQ68u/jKicfCluekRIF5Phg6bkeKULeWKj+AdojXOrnRhOQOgIA6A4Ducn
q1t4EYitwn4Dr2FlYMiVIVEjV3TUTkcSuAG+9wICvFsenLQjD7A3KOzO7tycHBNT0nwFCvQBDUYx
LHop5+T6dbakgEWFlMHY8qmsIeIblaQJTQxUN801a7XEMm3kesrTOoMI1NCqLUCIUp+1ENJQeGQo
rVGsmoZcLkctOKXXHA1HQJqlK30bx6HqUAr/BmsZzZPDCGn5AP6ML9dBmGsVuYPQz1uM4Ds/9Spm
kVbRB6yDrP42P0If+qd5ne30qMnRqMwLnoj04+5Dttp8iPFvQiKV4dqTvuy9VV3XlwY2sRoj+Iw+
xaMUnc7IXlsegb3utOXSz0XmM/KLNiEfdGW2IoXB0JjtsfJ397yska6YIcUl6fiRqd8J6PnSvT4h
AnywBzz2ni/sPe7Z3UCZGYT8ArRg9Rn3b6rYFSF7mn7xKXiVhbLtEvQp1NeHR9BmF2ku5tSs6Q9X
QUFSxQVLaeArmfUEht4yTgfx60J69gRMLDcFVt7R6GS5DJBb+1oprb0+nvFJ+tcZzMvG3Eq0bPBa
p+28E2FUJmQu6jCsni0FcUp1fqYgRUQKr/+Jud9OYUbriJJIHypNZTaSBOhf48pA7l8n7CRrAjDd
R99XdKV8iekXYn8/NFx+z9A/01fRODrjr5u2ucj/zzaQ7RLGw8SaDN0+42xFhSlelQKrc+5W4lTc
kdEOsPLTMoUI0TIpdUsD+veXrxeGn4frOJpuE7Z9BS+Ecpb37HA+0BoddUJF7zfKlN/0/ovZ+Q9Z
fpCOPAcYVXGTybOr6WHlZbusKGzMYl9MET0fJJdPK/22jVx4t1LfEIvW11NZPgk1dY8VQ5PSj9Av
+QfK/WwPIAyU02wGhutBhnJ6qd632dkhPy2cXxEt9R97Y7PlAFX3NG+ulPojfliScyL6whfYlG7z
SKtUBXvqDeenF+AoaqamdO5KCYClNzl06/T3Hf5Br6BaQZxG9SB2iE3EZZBZPoaAbd2muYesHyxm
ReILshCubHj3kvSBk/HLhafe35UqgZ4nGfe9G9tza3pXBoL5/u3rm/l1g9nDrEDNn/tR0KHBjYw6
33agGtbb7dhQdGrvln4uOyily0jMO7NNEIaffRqq8DUAIeMTERenNInpjSXB9lJgAvFtQNCcMbGM
LkOOmVYkP38OXQeqt7EHmXZ3JT9z2AYVF5FwecY/3VDFoDjBeJechgKTvxdeKKXQEkwkLRsICpqN
6tGuV30ZKQS3POfxiFE1C6PvQ7V28+wpwrbvDD/mEOD7TKZSqYkeSs4mat+YkapcUGug+pqpbYlB
TTa9h3RCbP5pXJJiXPt8cVthUvkP71IbP67cN+3KxEMa+eDfGD7/amQoWJ4Cba2lOOJ6pzv89Mdz
5TZW+vzCOW4CJrgWxfybx/hD5ptmP2+hIw4qf/vhlVwb2btt1C51q4fenFOsxEyn0/9qinmYSGA2
kXMSgegPZwf1rwPW6ZeoYPaXp8cgFyGnAF3W/pvfBVEFu/wGT03W270GIcobSnlpZWzW1Ire0ApZ
Ufq4tzJIY3Xk92yDnMJxa2nDWHiEOAqh0c7T5OEVVwcVhJsIiCcwAFukPkQlPKfiiRXgXWw+1aA5
jQLp6RZjaatNNNJLhwdcTtrOtnG9X5AxPGSPBXW2DvWpBCJwhWEXbRNAiqN2NGcF1r8k8flP0vJ/
IbK0blNVjG4oxRN7VvO0OyHJzJ55P67iY/VvtEy11qFj1VnlUrPIfu6Ze3ACnRc+UUcCvuyUFiNt
snt/HODizodgwmRbLO8JFILjI7UO65ITHVUD/TAEcLDcOLTUfNuwr2AIsX+wPDBw2TFaz02kCxev
3AYitBk5yqdNB2T/+fL2TD886L/GnSCwYolaZQfzTCvfPE++13S0jAd1d7KYCZGwlr/+KDNQMH7z
DZKc5zdd7RlLBfHzP4EJogQb/cH7Ogmm1mfyRtuWoDR8Kn6mILZopuqefZSfeoeWp2JJ5CoZiPfJ
xRotZ4+0AvK8k03nyNJHRc/c+lrqgORifmJA/gMA3mNiswARSsf28QhaWvoRBdkxcq0DJe9ge2qn
MNUYqjUC29Fl/0xvaOi+UV052bHqOu4qUnznBzW4+LZwiOaJEI3bfQpVw+sAAjbLZ79phG9rclU8
3aPaoU4Ml3s0BASchrJDdi9vRhDQBYa3W5mdUOqZgTHb6CL0HmhmfvpoZIaJOt+yR6Eh2lLC51Ks
AWOvfmoVREarEYu19U6VG3qCv2BGRV21tg2LYUgGeV50zqLzdykF7Pk5CtDgcsD3XUjAkkIt535k
0ESgWzPnEkHOCRHNgeM1mWet948B1NmPeLdHfWvABtrjrHyB14Ml9CcVzJbVrTsi1Y0sC61ytpmo
19SSDWEcZLr2Dau7ds1t7gLBWkP0G6uaqh7Y7YIzmLDonZJoAhpsyM6QgT8gvbLpfXgswcG4h5H1
huNHG0DpOPQ1vsaOrsWuPytvMUNQnAnYcnMjaI9emFCa9xL/oOaCrJuHR20PVJItGTfz9lFWKlsE
1DB7p0Y9TzfYEzaEdtLByVlwG0IPD6VEDuVzPlBhJbDxuIp8iWuzKUnlTNGkZAisxYYGCK9uHrMR
vljWOVsO2iuobIzKsWvolEjJ6rysPnpIaqKdb7jg0pi0a6QVZ75phFus4/UXuekYPCIknXl1x9Iz
XDlVmvu6MfetHt5rBu9CneZB3OyYSXejardhO89p4/Y/vnAShrX/W+Wa3tZdeKJ4MtM8spt0HnSP
yMGnVQ+feNvx8tlYtcyc78ZwN30feTI+xkuQfUxO31afrxKh42R2K2hstujjLVinhVQTkjXR2Iz3
wtseWz5m4Jq8ZQ7a4oBbLGZn+S/9oJolXpTVhHrjyCFeiZ5JCuYhwoJSk2nM574hgPknc0WA2fe/
nCXEKWBe7tX4bX8LM1YR/ChbNv8ZyCXn/8jXN19J2Exy/oU3DkiolNjQnz8uWa4PAYC220SxnXsS
AVdBCZ20IQnfpB7Lnjf4SjhXFBieC11MCipBU4cbcQ8VYW9czQLM70SO1SBLUcmgd5NS1fJzcLRb
Qoj7dnad7eiioqbKW9KlCtMp4hAS1kup4G1RNOS5HXq47HRz0kzQLZjc4Ef9m7elaSYAoWU5CQhz
PhuQj+yDX6kqUYAWjy6q/w4KRImXRYJGMrEjVJ8QO82b5eETyHWh4MVTc0i1hmL2xNQfmUdJ0VLd
vzzKXSFmbRxVATrSp4po2FCrjXYgE7lZKrQiG6cFM/1xnOEiEUgj5EGHAHU04+ljrabtcNq3T1dg
qHjmbtp1G3FCI7GQw7/zlFpRBBAHAX3z6AgHm/DZwkMkjuW0bISgJmnVb4wzUQq5HnZJoBzR149I
+Owf7aTXWITGPCdxy9yw73I90R9gF+mlAJEXPUvL8jkg5t2VHSUPoB+KWbhScZESrPKbrHdfU3VL
HTPavRRSKAVw6PvtMRlRku83AzEN3HwDBAbls5fKiuS8sgTkw+kBga1OVqolRz9CuXugiJAzeC5Q
hCr/syvS90IvzjW3Jh0+yfB41PUMyjDQ7xivaJXsYVCtqbFLCBynCwJ7qFFY8mD5pwT7AMmzkzWd
j5GDIj0vVVsKEP5V+2uuyCPKdbKifDUyxw1l67j2+/BK8YMY5+VLBQ0MjoQgPkItcQwi3YWLjBfA
7H9TDL7phMveO80JsgdKGfoS1B+gP1r48vlFQk0rzcDuF9S1obnTZNwD/V1LlEYdaijR8+sxnmHo
q9v6prmifmZ5oafzpqn+yyyQJq0qSMm4pA807TSoqnZ1JzSB87GeF5lGAnajS0olVOBPjeGxIBaQ
fwEylDudX9DnBkrflsBTCwZKubhf6G2vh/G/bUU2oM7fj8NfgfzXhjsCIBqUzFOf57IdwdH6ua9i
ydT0RIqpm86bNJ48uDGFAli/CSQvyUEbBk3Z5SYDZ5JWyGamCpev4zzUBifn07aMW7xGTUPL7X0d
f4ClYx1rwJzSDy6AYg8yPTRVDwZTLcYHjP/udHqk2psPwaAnCVwkE+x+l2dDxLH1DXUYQtSAacMF
zo4Df7Ckn1dd6tQuWgUFofMQemHWESp50+cjyVoG7dQca4D3uLkt5updbZ0abP4p7KC18eeTma1M
vbl6lUxm5E5shHIvkXcoSo/m5Lwg3oo5qUHjkovtsrZ3XLvYwH24CcEAxicNTydhnJW/uQ8pkEBM
bUO0HxfDHUYQGmWbF7hBTVoRRhgSN457n9iwWhSqu35BeP67GfyjNYZ4OrY42qWP/uFwdefKW7XR
YvM8s9DTw2RjEb5Nziv5q5hecg9fOh81kdkey+dZXitzro4lSi11YcbcksRgOr/cVF3Ux4tf3aoU
D0swAgZSeRWeokVA7m6IOhgfYsVhTIsAWvP0Ob6ivDs+nELFOP7UlasAmMzt5A9KrSbKJV4lTYU8
f6jYFV98q+nNoMD9nHNzPfZ8FNp9dhX/tBERu8DJ98cBmmZ3Chj/0p6g5WtE8vGrrd3qqi9I3IDf
1J4K6ZRS1PZe7lEid3Q8EzUoBVTD1d/F1n7N4gfGwT3qx3KZQwUpRmwh/0V2+0+P3DMg/hjNQYXS
IreWBGsEvGmavzRLLHaCT5sHRhZo1jMnzezA6urm8pv5j5JXP4tLNWpT21ehwM65tx8oX9hdSZVr
zcFq1Wzn5ESyDRw1jrcm0VSmedl9fhZDQTE0M1uROK6JM550y8y+z9iUNKwfd+7P7rFFlWN2SIAI
nq7s0GafWIugBOLN9RENeMNttx/Yh0UZRfB6ZU+sJdxbRlFGHl9+PNDjm32iwMh/ThVb7DZZqyhg
/dQOn4etJW0fX14/mQCxABb7MYOzsiIZ6nCTdRQUKziGbtwuO8+0pcR3PgPCw++dhq663ismIuNg
0+a/7a/1uWgZiNboTNh5agoTZ/ng71sQnhcHHyNcXVoN6pcjBCRXDftaINh2Z7LRuRb7zRag6vaJ
1wx31bnLQycc1NfegfLGmzZobV6+Z+NC4jCBLZiJOi7huy2B1cJtmHi/tYeF030RJLZhmvYBQ/O+
cbkw45D0Dg7k3SHQvvG9S9iy3+dsriWNm0yHdo9ToMrd0fRSbRaJ2UwFzCaWUC1YI0nyqQdcw3RN
3w5apL3ievnOWe4byaOumZW7Zf7aob+o9zRxGqUv7I/xP0NCEyOk4TASbDkBbNw2G0xJmBuOE8tT
VzfMyZVZR9b2cB4NJtiNdrjiRQQk5MEcTrvG2F0OBuAPmWwrDHVN+ZtER0mgeUZMzWG/H255csQo
wU52ceTo83ZMRx6z4brXdn9Tzw0HPw1qVgUzztrNIHrYfMVoVRQENTIKq4H4i62gKajVxOVytkV5
vpN5ww6+HPkFa81nsTsYZKX6KIMAq2mfK/Fdf8dD9lUl2DXNUfkeJgwvpjK49n6VEpC6bE90zhT2
P1ZOLeoE13JvBwyOQJMMFvrQxr2jFFZiMZvuCIUfnKfLj8PH5dv8VH/xHe7mOCuiHgHZ5ElNSqMA
fJ8n06J3c1MpFiGRgei9+FDrS6TsKmilAF+xW2Qn9PHyE2URynJI7TpgsYjs+ppUXMLAs/7c13ra
f4mzrqOrI0V+lMHAUVg+BQqTLJzdbueOxECFJ5fYsFRZ8CL5qsobxoXQk+UfUHF6ciaEQ0R+IYsD
yIklFF5b0p//PBy6VeHGiti5cJ0TjElMpwYoqWxaVC1Svf96lhCcLHvsZtF1Rr8cYuZeJIq57pIQ
GqdGRJCxvWkCXPs2QpoOEcjdqNiT/3pVwnXGf8mibtbuCY4jnQuqvCbfPi8uIpOETv6ZtXoWTl4u
rV4khRLfZHI0ZW4OPNz4NCtOnszSHCRq9K6ZoTng0xbMd6J7Vy3XMT8kKvoiPXak8LVNJA8Wq/JF
NLfr5kZzoPAIKdvYgtnaQ3tTl53kCQ9OITBH8OA9oyinestGXiMzh04Ob4Rna5O9VOPjdZGBPfzy
qJVq0YcULDby0HKoWeRJNLRK6mK3adS7qIFRgN6acLkWTGkKpwrOGKfTi3AIL0NmBPSSMH7/xs6D
/tYqlzpivl42Hg6bY7wbL6CTlI3y7xscST8ltiFFni85Al6d3ZKhkog7z2eGzhry3lhi997uK2RR
6DtxwifZQ3VK8HBidsNzShcn/vKrgvI3FZV5PsDaIiqdPuFX4huaOM7rU7uO+zF29EvxO/P4VA9V
FjldBEfsaG1yRsTWTxy9GIQG0dElFcln75wKKNhXdbqtbk+H9Dh4PKZfXAGSUlA1W7gcZq+wuPTQ
jmuFuTTETYfvR09k17UImNeM55JqMfDJnG6aT4E2OyMPeDnkD78sWA8oUcxKKhkl0mezGSCecjfN
Oxf6+G+G6Dm1ENSx1zgTUEZ0TB97Vtau8iPkn7gXh88WZ3GKPzti8JcrAiMXagbPo9tQ4+4IUgr5
tLXjVVJqgdczl4z19sc1hcp2/oq0pCStHBzW2LHPRCKPcR4QV2i6M8I1S/ChO2HNadOUb03oI4Ia
l0/yEYaKbLtjQo/+a0znkFjUZnLxF0tHSN/4OWN1Pz/oxyqVDE/b6s5j9SgZofEhNut9G6PqbkaA
N+8FAyU3zqF3idDRP/PhLq5XWmgLYELF6kDYHBIGgSgPsoESzO98n8QhYrm2Y4b1Df1XrfD30r7R
xssmu5XZVGh8PPVZtOkx8rUkY6yDRhYhxC+ZRYEtt/gPgF/R59/EQzHfgRj3ou1LCSVatS6P9ih9
xP11NLDnBUZXYHIHOVdHYQ+0AuvQJiH9Zzo6oZnvEnJ5IP0YW/PCj158SeMhkxxnFbNZNTWWoicv
QueeCiKXrdgtQPBb1JY1N/mt67I63haTrFZH+9uLSZJfbhTa+NmlVm3EvC7HxSw7JgsubYIy6KA6
Rbbv+8dpEFxxJxEiXgQr/o1iyvWuPdwry6XWuaEI4IbHLGSdN6PylV712ENTlJ7LcIK7m46oFttq
3BbjsJSS/IWziNrOnwq5bFd+oVNvYmbpdxl7aZNnQXvileuqvO3m+7TRBOIuqTQx/bZjOMUzPtlM
4WwLab8Mu3QVd60u9si/GRGxufSzrVCHCvFZm7/0HMPvDQ0SpX3wS8kKjptGQXOXs2FgC0w3Dmpk
5GwNe2uIIs6T9+z4V58oexIAMFR3vNQQQJBIU4rl3ZB8DR5z5WKROg2pvKOGqi3jy9S3ZeCu/Mb4
HaxhlkrS0F0v906rWp5FahZZTD3hxOx+JF+w1B7f/XV8TW4rqlYXcp6ImL+ZuAsLiBVywt/Vist+
Mzsrq8oL6TeUuMFlA/t3xEZS5rSFEo74O7vQI6Ilm1PW54Eu93Bg6kspMJMj8RsqRCIzIViVDldB
EYhb3EOmBh/Hn5Z/Cpc39yi2CUBvMsrl8LQJounZmb0JBdpQU/A/9PZrmIUmNcHzaortKedhRIg1
UW6rGYoic+PzqhhO2Gy7lqs3VAUoxMytLOGMC4OSfUk2dRzhy9d4aT1bGbwmmsXODETNoaDbqTTs
73a2lUkbIMFfokh3brcxEJTCULewGTLjR85YUvFlLo1AW6BFu76Hpsl3GYmsnip3DyeGwsmSSLID
+Go3mEJAe9S0V7hoO8D3p7XJqqx8p9HKfZDDhpISdPp6c2yW34B6QBzWqEw1sXBhTV7TQIFI9B4+
Kc4yoA3JFJ7cvSAzccUwEDLLkVzUnyZnUrld1tkDERlDeCIU5MBE0rRJcB7cB5s1O+K5qu3FyHhS
gQUcUsfOPgDEY6cuGQ1TQ/3Bd1et4DXTk6A31ifddf4D2g3HzoCixHOP/HW7Z3TiFojvrEHSuLOK
YnBn2k5Omj16Wohu/e1GRGjmduk7W6XLom4rUIZE8uLfYEFbJ2Wkg1ZlIDD1j39eQFAA86lo8Cmr
8frVrOQE3ge4off6zH6Fn/xdLEeNEazuJJUWvWm7qWOUTlSNuFZIn4TcY7TxlGfT5YClx0IcilFx
GHiC/6tBRUSH2eVG9IUAcsdrhOtMjS5l6IL+P7hAR/RtTTvS3TrlBa6cMLnX4GUy4RB4VbQTZh/N
gE3TR9GKCApAHRsG1rTTLcq9nlCsafgH3qyt+iIpvtYyxx59aEct2AgRW6rubHrVJmV1X+bW7Gbj
5NSdz5v1ULqVetP0P0ZmKekCwQXIrYY6nfkc/KlD0cy6M8ewAFtMZJ+KcSHUYu/Y+diqpKZmH5Kp
nbX6Bgu1rcb6onw+7dDicEIUAue+ggQeNqUjDcX9MW0xfBkiXhdVtnLSL3bJ5DPcVHryzAtN1E/N
foAg9P9PJmRr0d7qcOJCWUjrQEM92KVanAldsb0FhphwxdiuJAw32llgRjOCBS6KW9X9FdzKveLM
yCojLR2iB0Lxq7quNKcxKH7uAzIZQmyHbR1e0DXnMdVFvFJEP3Ij/wQzu/w2Kmgy7UfxdOCh5ZZq
gxKIwgal6YhtkgBPNxMZMOL0mjZI+2q1Z6W0IclqgolAQJzPf0KdCDhZyhpc02GxZEi+OgcAfMP4
wFGimqcduoUyc30sWxsiTM/2bHo4ZLzDCw3dcl4zhB0lv/bH7QzhsxPlncCIDReolKN74tPcY/av
+UViy/hvTUiSjDeQ8p+TtuFunvpJhF9vRpi8w+wiY5FJjZTVF7UhGuYsKghfunxeWjEc1qJEBk6R
ntMznhxrhgoqMRssSv5mWAvezmh6FEwAPqvSp4p+9osfo+iNk7d8XhSasVJc1No37KMTSjhgmULN
V6/F2QZROMQr0IKUeC/7g2K8w8sO2zp3dcm6nTbYBbBMpT3ibZbA1Q7W97UyL9sFSijeac/IeQc6
+jZ+klRzf4N4seOMeMTthH84TvP13PG/aS/47NylzPlputtMI4Dt9kf8BeZF0Nv4qZvR2z51msoI
etnrHpYGfL5qzw/QiJ9lfJU5az6mAW0zjHyAxf9Q9QC2pzglRSRDKnadxGUq+ygyakHs8SPwiSak
95Yu0gTxhI6KHHxtXaPmrLwSwuH99xtmNOifdS6PM2UEpUyL7o5mSzncdpVpFP01kWGoYP54Z+jj
NKy2kvm0tlyr5lt6sSvlEzr76nTkJnQcbbsaP6EYvJd6IQiVy7sHVRDAezHmdDh8FoH9ozACJHiR
NaHPuK4KoE4XKbNy6BvKQTJLt5tNOL4XhK6sv4x6Dx2GNayDyrcUOGmzprVZbHU4OmIBVfcOiK8S
44n66pKQXkWr2qct6kOzwXh164cT/1ZRfevNyasR0rO64hKHMekzYEPKh14kGhWm07btLztX3qhW
Lwaf0V7l7h3cAWG3mnSEuP+EHQ+ikqE1Jx3aR7roqAgoFV9XgeSe87MuqoRsrEZhJeCNmxz2BlGU
j8AK0WYmjtjjFXXZNFpqzjaiR+FvXAhiY6NLuz7b+IZxeX/JDAkRunTK32mTBvpHi+tbDg5U1WZZ
L7GqS4SYsYPIriAxfMcqYr+4EBHhtHWyUHe3xWlQkLZeo2k5ERgaLEoP0Xe8gLfojI1TG1lpoxaT
olyYtq3R59ZfiiYigo4WIHnEgTOjFvfTMm3WGu7ymjUsduluN5kz2f1AfvH/r+OaJtEvK6jbpAmE
CV7S1WtwxrzlT95A90YUStZr7sFPTPUkJdadLXf67jUaQ+xiEn90whAbWO6P81aUjnwrZePnT+4O
52fW0LOJ8umYTxKPwHsi95bNDPPAJylOI0CmzluvSePMi1lyyytX3ioDpDNc8hxnLjvBjjUlc45t
3c0AuoPKWtm7vkWtbC5iyIpMiQ/tKOoePe32vOpRwK0uaIkk+NjD3juckDQCHYZ7gbsrmnYaBJHp
H2BYs9G41Uupx1XapeIHwLrNvKHJUG4I4l0GsDKbavJH2dZisFU7v8ikj+jxRqo33KM0wIe7SX2S
MnkjUsWxcMyAm/u+doC0ZX5RZR/3s9FxGPJYdjftvviCjaXaa+3zCebAL+e6mhFbUgtrfHf3FuPP
zkfljd+WL6YT2825zUSm+2fgpCemQm3QPcoOazh0eg6ZxPaKTCCXnAVUH6HMnnfzyfOcmrzm1pjE
T1azZtRUZlkF4lWoQX65dHryc7GJT1O8pexGSDKUE9i4TH4t4xaBT9sFhu6hnYD83k/vQ/Dnrn2H
Nustl796YEc5X4+Y8nO1M/mdXZ5kDoeDoovOEwUtNuqDdLMwM9raJkUwxZx3hW2PE3hXIJo8xja2
E+0TdSSmSQsAt6yFYEBarIDWOTi+4m4QSYQl8Qnbfx6uYKks02UDAN0032lRRrMV8J3/SOA7CNdI
08xw8vQVdhvjqmAICwYI9qlRyAxc+9QFxIc50rGU/U/vHR2AFKPr88hSz4MyOaNYEXv+EDNXLoKl
LDWvHPLZ6Pv/yJp0Zh50UUYEkNyKkyAFiqAsBi5mY9NM7dL2+avZH/622Mx6aGDHcozNYThpvR8B
erpydfKT3NkVHEYiTXz9iDdqPVLGXBndpnSrgN8YE7HcaUS+SLTDg/0xXfrmLPydvTs8TlySXtxL
ck+JypBenoezuHvf1SQoE/bAsy/Gfpfh3f8Eu6SEL296VnLw654b392UT6lKRr2Mn9o/UhlLiYJZ
37mwd/CkOH8KXMoqAAUYPDhvXdu6hLzD4tllRJtnIjKmiBpG5+kZD6bqpV7DhHYZ2BiretjiKrDs
Jfku30AhJIaPiZqnD0d08zj0QUyclVcC9KR9SZmAbLwH90fVZTsIxFo0JZhLw6lqn2GI1NCYKypU
1zpl7bHSikVefjy1Xv7w37xvHZRe7kwi4Blk1Ik2lN6XI80dwAk+r4yJy2sXUZ0LAHANRv2YKmfs
lCTrG+xJc4GsS8AZF6DQGCK/HevM2JxPbmBah4gG7qLG0nLH4DUjfR7sBV6our1PNIek4LQc7GhN
I97jPdmffyGdUmKjdZVlRFaKwYAyjJaRB9JOWQXwgo4jUZ1lhE67BehsEjlK5uHlW2HdaVyvLlv/
R/MRI/6NywbDNvgvuy71CIaUsLOB8XQmMVxW5hEVxQupGDr8FDW02HMsSScptSZQWKfGl1r5yWMU
PkVG3cEKgwU0AKLmX8Te8GKav7tseAZtBYwT12yevu8rEaGbp7Mk4/iUKDseaGynohKxfqkFSt+K
B7zdalm/bfgMIX9pYZOSBXpXN0ZrNVTlgKvLdbrzGjHN5YO8ny0b1hKzTxVxYKFEr+LnPtRTDsvY
+Hm5oGmPs/mpevokJdOk1L2nxAuFT/tIKubGVU3L9sSgoQDYLFSDrhLcUVVVhffR/meIFVxOnXAK
QJBmoyyd1pwgY9+R37b0PzkiWmXWBh8PwJgk1C3V3Jv5yxADlgZAQ/PssSjUktNamM+ByznY3B9m
osmjJv8BLJVecXjTmStorDiLEXhQfpd+i8Nw7dDQ37Ma46XCi9WvLXg2nuTLt2jc5JkPa5nf56D4
fiBrhwivIIfAiPpNHeRwnhLY4a+BG1aL5UhHKd43I7R+inSTwzZfGMpOMxtEGrX9ZdG+20ZbMNfV
fviMn6LycrhBo8mIDyqIzys62oEqQCHQN4eTxhL6SeKSIPlnySJSIXZq+ruzy9PC6q6xOs16z+6F
14AHuLguW6b5mHJe6zWEmYHlcqdQ14WU1gwiDY2VAGqgpi8vxSHJ2hFF5508JoHDqldtXT/ebExA
thypWrnyXrBwYE+Mhdi6I20ey3iKCscovgdHSUa979EhfbihbvNhHKEvwS2nAV7ud7gmB24yosWI
U1kZMX6DsW1v+1VmoMJWKJc5dajLnYa59QPgTJ2/9N/+Fj6dN/XYf3hAKmZSSLNqM4onjjWgILDg
wP1rmM6/v+TqALsonl1MvNLViNfq2iwelohznAZONgq2xVzJ12U+1PgR214hpUe2Z92s4VqnxYhT
gc07RPoDLAkQp25FdiYfBDhAC1vcsWmHBSyCrpvtmD67JPhvxsXxBWACd6UZmHyjiQ6SuL4tlrBb
yVwUYqTwYKMDdsBTIXI/6lFGrZhcErKfWCpqF72WsqaMCtHEd59bnPjc0MS4zpAisXPzv37KIY4r
F9kn3FnJCU6LYYLDQzOqKNihIzW046JtPTq9kTpa0uQfAqcyX6OppT82pzENlaflC7hfmWjSvK3V
TDBFVavIxtarJ8uB2t53eytbaWPeXXI0+os2zA3ohY7y0+b6mHugN1NKtP4zkhz6hGtVbopkoxHu
8MWgtVu6eybGQkEWG7OqUctGDnIZ5/Nu15Guiaqp/noGIKhgvKYBSg98//5A//d7dQ27tsvpdp1s
V4gOY3JG7icGzAiG71eFT7f0OrJd2hCgRKf1S32obryNfmUkM9HAR3oGFGe0IP6gVg71ZykE2X0P
RTIRUvIiElZ3yhkMqSxpiq5c7xgqYkMTIBszmJhqd9EYUByHI6VU7bGr8F382MdfAsh8xScLYWBg
/D/dH2133JJ7bKa13mkH+BWLqeEOQzT+9O2X4kqG2gllKpx2kmx1YgKMoUrO8KHZ8Ah1daymZqST
+Mg+psILgc4u567ehTeczz1lkjplxsr65IKwIkwDZFvcnTOe4LNCriTddP8K0xkzLwcywjS/vPD3
Qryyh+xCZoO0Pb7gYKTxVaM0LnfWJoub2PZpet3IWmZfmWssKlVXZNxOREISoprknPNWQ/0/2Zq7
fIQmPQkQNjvAYkZCC7ua7Ypl/Fqj+scIna/Bna+7xJASykuHlFzdcyBj/uoQDfpHvx+o6eetINm9
2lw5ttFJ9CABKv77FwoZHiOdENRzKLpFXNvnztyRz4IFNS3Rkc2c0bhZKSfmQBiY4qQsHe4MMfwt
cszuu0G1DwMQK/gyP5xZeyqZpk5quWK7nocPcyMjJbozjEwuHZtPVaTmQZIrE9o0lnVumZifVOhb
WgB6MnpUSX6YSYGMnSuT4cdIXQFRuwwQloP1emseowHubAY469fh/3djL6Yf4DQyinwr30ypn8vk
X1jIAu+bjFsVQqzbRgu6+Ne1uek6AIiiC06YzgL0cqEPa3yH3V49SMVP1RaSJ6vTO2mZOk1PulMp
kyZePu48D942E7R7h3x1pTl8W+gr4c6QW2q1CtMFJvmMlIsbaLN1Mn6EjclbzvujIshwCPhGzXP7
jCBx57Ys6j6eWpJ+S1C3dsE9Jw7kMFyNH8MgiCXmZiw59xpfCU/3sMhcGl5YkH/LShTQpXKlCu5c
K2FmPu8o45wCDF9YmsDXRI1oiR/QHbUw3ksnWHABxgWibIFGkcCXtWEvpZ6k4C4S8pBVunIqo0ct
YYKZcTTp1plyz++LSnB1iORwhqYRH9m4OYvwlS+0va1mmKJww9kxZ/vkAEK2yxh6CsDyxh0HLZgg
8UgEg9Ba8ElA+5mG0G5C0qMFKqzgUkXX/Nxl5TsUdwivmtJluSllbkeQ/qyrurhD9rE3KtTBqJh2
uL643mmeBkm20kmDP23WpUrwBMggTk9+abG93Z12cNzGfTX6E0O7cqie58XmARVe+uM5zIM/wWxs
mNxGiDQYfwkRqaUIUdfJaUpNQnCa47XjlLw9Jpikapub2wY941h/QKWx73t6wBIWpsRCDDQnTCLZ
YOEFk+pxcD7LiWJnZEcEBR0Y1KJFVOy7HnNkvy6JUipcqdmAjwV4ywn551vfXhsD1PIoXDFf9dEa
iysF1YwZ+kxvZ5TKrTFdkWFI2ikGi/XTzwVzeEiVUQ9detsv0u+XDm4hn5z2i5eqqO+hVKXdxjS8
xcCLUnOOcApsga5xGYG7OzQasynWV5A3XXOhg0mYf8hZpgFEKbtvw4qC4mC0RPJXivMNMKCJ80Uh
K1XSFeqZ94NGKWQ4wFqpVD3GCS2q9FGy2qoS0cN/k7gC/HwIcEu5odbV1vuM795EEA/ws0UXNctR
y2YbrakYsCK3wUsLw3qWBmL9AoJBGjxwvTyYTMA5/460Q4sOpaIQJSofcWiqP6DmkYhdomMl5WFe
7MVzw8I2rAFbn+JjmdBo9EzVeEeirR7G70Tzd+f58wNHedREUL8u66JWGJPl+ofjg4yLs2v39cpQ
/zkYMBmG9/OcokBbC7yC/y7Gzfr3DocXvFPWfYSeLSWEtN99k3jl3ksWkjo0OWaqR90PmVj/1zVe
nzm+YHJYmUTGRhuM+bRFMt0ZCvAlnk/0CMeaNVho/OwpqDWc7wM3ScZp7i3D6qD1eIlqmhbJwVNn
QAulBDN1miilA3chwA9uftrQxzwBQgOKWuaSb7jGvupopscUowjIWERGv11GApE6WP8lLGoSTH1V
ZXq1qVqeZVOll6qEHj8fWO59gGxOJKx7sa3tp0fBu1G3wApyIzL3JK61hp0H2w7LeaZvtR9kPpQC
XhETHc+tXZjigkaNwaysMFQyjkXzKk3q8C1SYbj6Tv7IaUrI3B9fIEmbjZrUQ3TDSybzu85JP3mi
JFmtHJp/fqGO2I1YTGP/RUrF+3yZERibAs4llgeMZ0+BazYCDgBjZTy+zQHguy8IcI9izQqJ0AQl
vRKl788JdM3OfLaYzATrO+6ybnkoCLOWGv4an78TrZ5nPKQ+UXLivTdbo6t72trLCqFI4C7NZ7Oe
iyVRmr6ykXuLB0CO5bn6pS68kMKopiGTS2ZN20d86Iru1RaI9nCrSGtV7t7397+lcPgca8v20hRW
gD5QjDqliiyvS35e3Bj6rrKY7XjxQWDOxdlaORqBbSsHrndhjudF87xt5fdv+A2i/s8+xNLKOqSP
p+0TpB/XYfzqW5kZYsPC2cHi7LNYZv9xKJ33pdmCXR0k1c4+LBI3hq625Z97c29npFVPFBPvOsb/
NNv3tshinmZ7ZkDTGT7brTqZG5JUOyc4g9/VsNZAoyMZgGjNy/Ha7YtU+eFC/E1+fKBhyW3ClDvF
t4caKhe3506au5CLkRrFGu9/36Chfsk/nme/QbtnHPGnxYgzP+5EQoHWFirQT4qQyuTdyWGxg8vV
LawVh0xmUbTK2lZfeUuDAkmt3eNINowB7+zzizYoK8hVzcgD7R7Hkq0wwSoqPhQCiLqzmSeNI5Wg
VYcEc3s8gb+jML4YJ7ABX/bRKW8x3tRMwlEkLgSH9jxM792Whb+wc+m26bYmkzcSeJaHlHI5fW3K
24x7EmGfIn35GgETwJujsEy8bNeA0dpe3JRjzSSqWgoLddFiafLT7u4gwEOxf3v7VBYdL2AlyZdt
y+ZbFG5m+uciGH+tTgAwOiYmRTeNb5wIH+IL5bV2QOc92+zgCoJE2oj/2xrfXpVaIEPsRYa5xr55
ZACYCaZRYbeRwJQFCZBmW78cTZ0rOvHCu6u5YC1VEfSeSZ6/dGqcqkWZW+MQG1gpxuaeqcyPuWen
4GTBy6VPozuNg/X1JRebJ+ZdJPL6elVXFn0MzpoPwVgnj1kf9x3BnM+aA1nb2nphRr6+x/ZdEHev
A5NVlGf7Cmu2JHKI4+QfLdCJQEJzB+jUY0QaJc8ltVj6Q3kSxjCUgjvek6e3CjQyrzSpg0Ua6Yuj
EkH5aDV0e5fBiLqKLhVBYSf2rqTTRP3I9Fw8JmnFnH2YBm606Dha0n71IwgIFXf/jEEL922buBPh
N5iQnxQ4MKK5yRILZbEAih+hEjJci8At0u4xBesuqMmPQFO3PBy0jlnvWbEvG650zZfLgZXXZuu4
acOWYd1c3Q3a8c6m0ERBTzTKPUZHhF3YxEE5Dh+YIghc/CDBXVkYDPwcOmvwBi/b9vPiHlyoOfTA
zOvvlNtbOQj9xvGWEBSc8oDkpasSn5J5zBWITy3rOko9Fq306spZWwFkhwPqAb/jtfeBtWCqZxhA
7sOU1tbHnJTFSFSWt9DYx8V1ajQZ6YL6UlgruW4CTTu/h0SrKFoxbGDGQ1/heCXT2eW3zTQ2eIS+
oeBacTDAZdFGRTB0IEHdt5kym81gI1EmNz0Qyo1cDpqjsi8h+KLN4/oEnKZeL0dbVmDeVUSMHLQx
TVJGZ+d9bSqu1j5ultf8DnbEunvxS8tW3K+HVm9daN6Z1HBsBRU2QALkPafoRnKA21w+Vd4A4abg
2Mh8SKCDd9l++1Uh2uXbM7iVUx5VD1zkKiiekXBfdsNGRIi86j6QF/tfPYxSzqrsXYLqdtieJH5L
qHo7TyyBN5LEhVzkDQK9m5GiWRnyn3LAKqB82j6T5SX7m11LjfFnAB6X8oRK65oTzcG/JTWKZyMW
T3IL8ZyoY5jSJx4GbpoyhxJAgdXHYumEk/uWGZUvTeX457U5wPFKS0wgIwHhknvFMSPE/kiM4Fwr
LmRrzBTMeUGJ+uY6Loyac+ae08WgxAgKu/8u3Lxx8iQYblCA5Hcd8N3v68xUg7jhAAJxOqmkCxp8
0w0v3MmEyWMipz9jh8S185ph9Xo6aEmnGOHnQH2OXyunmQlggiRWr2HmhAG+ZwKboAho2SF+QJgS
YFxRILr5BPJ+FnM/Zlu0GNdzyO1Timn+oCYjrm5/bbqkeOZVnuFW800I9hONPorxqKqOfNFCtUPB
F+vZ0Rmjq/mYssVECCA8a58yWD2gbxFkl8cWFCCwEcBn9KlfSc7oXC+KpQono/b9osZ1qKcE01E8
6hfcAeRru/fy1JUFt8ey6vyaK6nHMnYe64CNPJAvCNwkwy20Ux/ZYWAYF1/OEJQgboa9GW2mOvqs
qHht64pjgHnbcgTNI7uRiY4AecE/pTNngbHJbdkkzF05V3mGjoUq0HNzaaYmAiSP960EvopUpPgi
b5OoAJsaPTW+sZ7gepXoCLzBEV35DrTD6+0ARDQtNJUaPKeapO30neARCM1wlpqbRwQmiKvtk02g
MQjZQS5BGBh2z1lMvKrKKCHLHmqTWafz+NhvnKzFErV7UV2nlEhq5wazcqfEBxcc6+q2YR7hphAr
I6RfuD0qUurhJ0bDXAsHNcD+ZyONOT4Ka8X82j4DvOgIkmaf6uLItnP7AIoMGYAJ3mWZDVvQniwB
l3yUINWW4GwpDfyCGGgR4kRxyICIFREnVlPMIPBCxazGcEeelFEXIaJ3675PSNj6sVBIeBmSlr4T
i1rK4xqDy7wlt7SKFspNzNm0mWuv2ltizZnoYp+NT9cbUN1CtUJX93OpXDNyn2bQQ0pPPN6EnEtG
GHQmHphxjAbWvgAxBdis1sqBYnOkfH/9RWZXkvy1UkW2o4p9rdC/HEh06aoaES6pt5pQ2ArHkX9B
4tM3KhH12Uo2PXSFe9tiptyys+OSxyXqLYJIEmhDbXBValfdaUTxmuYEOzRkxsTpeqteCBbeyD/c
C7jQNSTpmwdD2fH8plGOqbh+vfjTaBgl0iZ2RR8d7lC5GFbEEWpYoAPVSHjj9wiVvdmFCudERRBp
g2MuISQgaXCNGt1w+krVpE1KpbHpOPPAVWjNjLgRsY2J846MsE57GkwhEhfA+T3A/Eb6AG+gwn3H
uNC9DY3eSEz+v0JPw/4ue4oddHY5TIs4MQ746evjlV4PWwmS3vay6wykQtMaTUQRW3NfyE4TnkfJ
CrPCMj8MeKZGhV0SK506Lu/5y6pDMjZQZLABNNVxGeGn38z/RG6QmWHdUAezA7NuS2GCg/oQDwSt
Scd2P7PCqkJ+0zxsAIBlj97VBf5voGdBm4C5Dgu1y09MXe+yr8TM2BK7wNvHo77SJijIVTUwP0/7
/qIkrsY1jY1zuoNqlOutiLFF1SlB6rHVFD42a5SKA6X71uKCSPgGT+5tc8YEH+thC6+8Zw3f4DII
BWQvSH/4NvS9nxKYr0NsjeWOkMdcAwKLsqcLlmbqoEUMEt8zYljbLmlqERDw1c5FkQuGoiquECSx
lOOnb/Xz0r/gPMs98KySTUL9raygGoDJVehloyGIn5VClxPmn3qRD5pRz1W/wLvpG4VbLyiJ+hCM
iVYkukac81jFaWMULXr+a1onn6KN94XSSbCr2uFXNe5zcTsfXBPpHZIbP1vsVBKOsjCwO0jEM4x2
NWZ58e4zKnyuV0R4sryzdbySdKipbSC0uOyF1ILaMcii+vj6ZzE/DdTCQXDpzFP+KiMCE0JQONXt
4Kaxd+aG1WqZw990KBFiPuY4CQtfhts0H66LQTQvlyjnh/Bz1yRdAIWX3druC388+BYqJoXlHinx
NUJ4dSNHDFnyYzjyCn7NE0jarnHZiTapJuE83Q+ECEEyArSWxUe1dS0BlsgurRFHJkLmvO59Cenj
oQDlzhyN9+pajJgfccWedUnNsZZ+ifnaMeTcf2gHnqp2tAZXC7veZofuB6a+SkNi9KsygmbkyYD0
KU+AQu+UiqTAmboWx2K1nenvxqzZz6PDAvR8TpCkcXXTXRNyigZKL7hnWw7WYKBQCfrqFslJr2WY
cH8ypbp/hP+lDSEIUjD2G2d+1BuNLXS1cpAi4ofvmUiZ/sTAmu6IRhieOiHeqKBXrzDKzZZ8GC0y
iS0lWkj7GiCEkc8Ia5/OhG8jOa7yBpkch3gagrbJfKL6Z6hJfFevl9/s4SjZFkChGe/ktT2RY6ur
YMcIjbWEQEY3ed98kQ5t7AjLxurIZdDmtwlDmJXmmlwr8PwtDtfnUlKLgr4qX3Hw8ZbA41FjJVd7
Pvf5DwmZgXthElUX/zwWPAccyBC/iv5BW9uJzgh6Mcw69LUE/1YxuXJsQQ4tbw6LskHoxaO53eeh
RLp52PiMiwSmfRR+90IkJNDz1mrvAVI2NGhRyY8f+lMyfPf9wJWUcSblg5xf5L8H5Oa+vufTupku
8ueN26LN9MUhyPZsUHIMf8soFzoZiRH/4Imf856hL1FYM4powjhwDdQXOcWLscE8AJ47D1K7JlVP
zxe2Wjrv10vq3OopLU/miusuTrxX61lq7pLOHllyvkFK44GAATPEiYVfRodRiFbXoEoFu6eSDj3k
TQK64kZ9yCbV0Txp/byrFCxlIQWSVJDZCJPk3F3k95JTYspSZtxg0vygpHnxLi0CM/irLJpRdgcw
B4nZREhQ/p7//e1LHqavEmhQCxlyr/fJBMK4P+nkwW3b5JXfhwLZVMjvpAvkqkYTunP06T6zJBii
I5hyda3J7uoSJZUWS1PrCXS/+AZ+rZ/YbZFGtpTF2L3PaYKaJlYuOehFuwu0/YKsZIGKE4wxHmwr
GtCQcLDkWFtx5Vy/KFXoWBJFmQRCBHiXiOVHYPzxgrbwPoykLXqsMY+WfRO27RaWH9tYWkYyA40+
nlgDSWxI8B6SV+aZXwg+6KgahB9ERRtAKz0fR6G7ArGco5L8fIHnJI6Hxs9jy1K+pGYjXJlbvZhx
0AZAjoeZDAQxRO99FZIc7SpcbLJqn0H8m40y3m6aXtILJiZTEap7SQdlgHknEt0CfVwnCAd0nPdx
9bwF6H08/fdqF6lvN4tASb2A5v83wbddkkE/grDwiPRNURI1x4uvToFd83tjNCyFOdmpkB2N9ISY
XcC8sednK8rmntfjTnOk0gvRxyxvxUfTA38GlAj8u2G8H9TFIu+1JxpVuGxMUJ0CM7kBooXjebGW
vKN3sYlXN1HcPmjGL9g+Cgd7HnGFHlgGmCffruVS2WPhuaooB8l8mpLZCNNZ0xjbPPd3AJl01y01
YXE5iihgqcCpBfOqrsr1zT5ioBEmxUwk5+f9SYWjre/AghgnznkZO6s2jg9dVqV12nrt3PnxASH0
zoQ/0N2fjR/a7VxYIvS9ko57cRmE+KIQ4WKVCgp0enq0sq4eNOuG/fO1n7tARTc3GRttoa6GNS+Y
4nQL8f89xPB0eYgKn/yGQRp4oMml4ldhxAdrUq6fZVXiOlQvPh/JrkxrFtFT+OjUucRVLrcXXU4Q
ngp1YbtvSpmGteYPf/aQ5uzw4FEQR0oC6pOVzqayNhUGrh3ZvVDVubhYAXcTsLj7SPqIHolLFugC
wyA6446Tvvj3lntmEOYz6kr7tFrnS2K/s+eBXj1RJ8luG1dgMMfyLdGtikFnTjAMDA0vAMUr2wgm
GaoqhLZS+HYx5Fqw0jrjV/VIzYgNGlbz91ZpFVLryiXniAvaBQme0PhUMdJhjeh09lKkKFKR+Hoe
p0wWnxQIEkGMi/TM2mdtQBf+A9H+2EDp0P3CxJUGFudmLDXjsiQWEM4sUDcFPUGWJlp7ZOxTuavH
3YmGrCDTg7upoBhE1sUuSFHKTJgZctmehugLztV8gVfeS9C45iREhlBCKYwN/RbJNnKCxzoTGZBc
RwVWKMpU/z/hIeDegVpiLDUfWrsXNVzJE9mvdyNXzyklRiehNm/21/wnTy9rRBLU8qs+JkxG8f70
c33nfzK7cLwwZ1AtcRSeRY/pD/cYU7oI28WfpRu6YUUI+7dRZz15EU51RyxPaPjwYLmwcnkTVKwD
otqgWzZZ15nXz7+r27pkTz8+sWDpyCnf3DQ4Zlt9tY4Oz76u+d/N6uW2YrAPVZwB1iEOlgzgj5/0
q7YCmjMEx1RjMEGVHhu3ylYOhtEEAj/omJ0sBN9vNeXw8vfP2fPV8Y6KAL7WGVBzza5OaQfYFB11
jighb/cpg5TumrAmi24tiUIiUopDKrgUPnsrQNTzqzd8fWOeWPAjoZMbe98YJbdIwD97cLbWYZPZ
M9sEW6G71SZnz+Pb6nSz/KEQX8ntsyNpjyMS01rHxDFVRXzuc7e3GpHNcVdFhkLg+KwF/LAY0Mpl
leO/whzf187KXG8f7ig1m5pS4hFWu/KuVsrXygnuuYxMfJ7N4tABOZeQQV1htp8EHcVXNW57mvwp
/x26HP9fmIqmmvCjOApmu3ltnwIpWZBlsKvk8MslYl8zgUWYdvDwB521Jo0vwKmEZnlDEqyycoPq
g9QJiL95X1Jhzu8xJxqGlF4z4Cb3GJkXXAfVuAiO5l/IbMVSWPYNBz1Jc66CY2ljYdvzD8tO3ILJ
4lrIBFt1pNzFVI+N85LC/hJiEaX54R76u/pwLUgKWNjGerWpeiYlbco2I/ZFZI73mmqpSDzAR08F
fKdfPTpA4EOobsGabdrA+9IQhmBxfH2Salgc2I7mmnQWCBtO2ZngU/OYHo4Euv93bOm3876PQoDn
hkCD9AkoptcWuRDxns0VjnKYFzqsdlFj5MUUBxfX/2tQyT5ExTaROkuFfbwHGa4J2Zgr+WZ5Ejnz
dWFZJNsgrOj7ROzbKEXAkWXU1+7LF/Hb0rRP6sGxUSt/iKdV2pFZ+dLMbbr1ve9gXiLn6GQOmxGE
2FPnu6TLOzVscas2IWdv1eWNPw7t7LofnRKs8I5fhBSBuINr4fYQKpnG2CirBkw+GUs8BYqMKBLn
scWlq0WRldR9b+ftaHwZjVuPdaVUZwGXUSvXBMnOrgMg3CjP5/qYSd6Ia/aCdaX2COhLZVrjkExY
wjFlS9HTph2XhdcKgLF4axzUcmKwdEz5e3Fs0WGzlQbE1aMDX2z433EXk5kR/CATg9GwOkXasvJK
TiI1dsW31dJGZKRWsqdzYzYrpkJzy7fwGwM2nqZWQX0EWXyo1LxJWzR3feNRLe1cuQDjIMvrIa8g
DLQ2vfbhltUoVCd/My6R4TdBGCKGV1irApMKzSsYKVYLljiBXy3lYRu0zTM03Ppa/pCEMiBeaPnL
i/fG/jGxDjAq9N/0YBooY/GBdY1kQJIJ7MhRatFNGd5QMiZjhiPX1Due3IEoMRaqEVQrSCCzskNu
N0z6aNCCOWwF+sMeM72Yov1ehr5L/3wx4X/oes+T1aEaFNU67lTAZ3ujMNlO1qmibEYQENcOXX+l
GgYPLgQJxTlPo90zW1SLTZxukkjDMLL/P6ka/7DxProiq2LsiXpcGJ/X6oWXW7ZmLxNFcjgU5+c5
mfdtUlW706TodgCLr94+mwOfeAxwTXCGY+hizSs0fOz6JlbpB7zUaTyWnY3/v0coxt+5gRIarLH5
pl+wkCtkynoXyJ3fh1GflWTeKsYwWUYP2tR/pPeB+/2kqVPtndMQ/Hgs7faOjmMF1yJN817gfSku
jMGkbqJFQRDxth5Iwfu5cieRBBOTXP0hvzPzXObBrBpdlgAb2foFPy6fKo4F2n2+emRfE2pK6Ps6
ottV6660H8mXVOhNx6C8bM6spCCIX3ijLn2aCqxLt5Vksce7neYrQ+yM7WE1b49Oa+bUDBfDVFwe
51/Zu4jFUEYtteFMp5cmkHjhhZki6rRYYGBi611Cm4vB4xpOEBYDGP0fuXatcauLYHsjzZGNCaWf
A8v6CXCc9Vhwf+2+034imYFPyOwmogLOIeHAKG+OaG+8GYV3MO3zJWC3/140XAdgirfpw57SlQVw
GZ7kDxR3boqQJH4/TEruqxSHXhUcLetTpgIHpemFbPHmvExAJ7gulQKMeZJgUVJ+9xtlTeV1ZuHt
vFGC0GC0Gv2LzrDhpr/H73wxMwVpxthaq1DTSCx5ZfqaGAOfgpl0m210saiEENHm8QdJ8iQy93cU
RgzHvY2dn/fYI0IFvMhd8dSoIe7WXmUwCK4Nkd2Aa4egiXpN7uPs3u4yyjb+tVnXDJC8JlxWF7UI
wUjHyhYgPPVOOUZIdgud/JPWNMWKRnFDdWYpxX2EzvX2Zn2YkKxnXOpZzBIsK/7dHTH5hFmsCcnX
izAxf9fhjR0Hs6gRiQo0IaNqwsUH5170TN69F5qdIX/lC/2Irf88pO0rhD3kGNs3V3qZF1I95CIP
EljuSk5nWzeuBTpiNRKv1cY02UqM8ymdhJUZOcJy6Njh8Oxbqd5BbZP1VXq9Kp63BBdFFeNF49B4
sPBUajJk/8JwJuyVVNDN8RWLBembuuPLtosYfzqsFITyEfCeu/MRRsiSau9MCde7e2VsDTBiCtsV
jWBCtPR65QDh89o6wgscfvfDDnsfyrJr1TbtTSSHetG20dWjuCzJY2AdD93kdKA6+8NKa3rD/ckH
LTmm+EOVhLDfqPfe+qj0NfVqxojGbdOo+fh4iKXCJsNOEkgmLs8VjKIUV7JUZuzDexoSB2xIqt+l
Tpw6kW1iL9Pv5dfyhIDKeP+hlPIdqkgfeVli+pAv5FNrdOY8BTUIOopBHNC7elCY+4E3fHRy13fy
pqO2S3UKHd+Jrx01HUbzhN43F+yjDAyI/IY4DqbRPvKIx2F0rxHHb/2H+g5feteN3PrAI9yU8B4t
kCUqPRKzwXhMVJX6Me20bS8etq9nqPDhW2XvEhhLkyxop9mmJwVrD/4gIxAoyFm73roZkteEusfL
jjYhSCAUAkTOmqS58eEqpWDKQlV8uIPfd+nxnUxXwtb0nLZPWzhd9GgVOFZ74XsBH1LyDNm2G7ga
CrJ9HL3SaDyHXucJ07vZLBSeq0UDYtJwaXHn8QzDqleNw9zsnNZzq10IEfVoBV3YD8ixtPM7NKhk
S9Jch1kbekzSPx0HQlBKpQb/CGkaf1agt0QunL5OssdVMOoYE6MIsMbkua1sCq/ct2rJPeG2/qbv
5PY/G1BVPnOIXqDs15pPyrNXoZ6Z8Pyo8TSsAovVF80xAsO7iwsSMkVHR8azTd75mUFTYxojOa8M
KtqfelyEfIdp2AqZwIkm1j437+DjX6B8ZMm8mwm3xN16eYPeaMISGtdLY60UmJtpYh7E8UIHPQbU
VQbZjNAnhk5SUovrO6vm9CcSXH6apA26Ik0J8hino+i5kzKYgHtdpV4OSU6piqsldPivy7EKDM6f
8lM29nOcwGMl28KS7cqiBHBmUUEoLgeFgZqGg1/Tn+rpxsv8fB+daX5AG8yWZyHNXum5QWpBGQps
deITSrMpWPHeoq3IU7a/FabfLqukF8Xhdm1FgfRqDyu5JZiy9YOfl75PapcqgGA+4AmHg+awGweb
JFn1ASy0t+c51xroDXT+x5yxgHPFNa0UNRCMD8s05eyIsG8ul3mQiw8x0N9JC1qyU/IDAvyyBGGl
CVoHpyzeZNJmYkc9QJG+JFZVL9LEEIY6nrygnFAyEiq0iSEoK0m8A+N9QRycEpCLAgnmExDma+TJ
4atKJV2AbTtlKKwKSRk4pN6ANh/YOLnpKzAxzfMKidVTVKnoJi+ZEY5wLavaRdfLYnizIpHs+BJw
3NAYWfm+Q/8tWhmpPnTH3rDv13ZRQcU4LHzGQeXXgDt+pNMTvLqYthmb3Y+R0wgonOsXG7L99iVM
Y3Gwf2splVNPhJkWPRMszgBLTmm1FcS842S6LWq9hrfZZNVcNXeAZ64jNiqJw0rCdGwc3IBSnYyy
lJgOt+P7pjhTWgP+Yj8u80hGUcp+27UvHW9O+GbyVEMMo4ku0VK4sKQ06vkvLCf8nZoCENooXMkx
h8ShBVhdTlB7FxBacD1GINDQ9Pg5WB4TP2g5lzv/D0r1fJzYFxHC1QqN/h6OndaDlyiYndxmjeuN
QlPVZL+f3GSkz5GoOOuVW2rpcwQ0Jp2o6s7clKmevqEKMWlucImz2JFNl09xf9IKKYAyvC0bS2/w
BEaU5DSqQMwhDxxktR6RZmlsn9ICGNZmNrfMo6ObsSqFQTD4oZiIKdYo9LJOCFZlim+cjYogkvz7
UV403XlVcRKynV/BikPw0/4tRIMkoL6Tf5lzvVbv7P8BtS3m6HN9STGeQ+flcdVMsCwyxRr9ihuR
88E+QYgfqbwVEciXONbkNjeITMqjTT4Be8XYt5ZrbfqfoLRpyg4fXOBGPvH+PzOCGmXrHMV1cvAK
zge5YencyAklDKnehVbHnMBhZ6S0PkRlYqsqA73Tj6hG46utel9iuTbGZNITjxqkStp9tqu9pTBS
hgAWAgiXf2yWouOmgLSPSlqFxi0aEOFGqhUYAgEg2OdGczreku++HYvxvQIv1gBQapTCtlJJ+c+6
JkSPtNQdKAGD6TQivw0QC44R3D0RAwJPUqtJAQ6Kh9pXUQa0qSOWkZC3PQnFDaYgkusCfL4m2P6H
vCNeMn/ll1GiLG3FDGtV/sOppz4C4LlYjf/DC2Rr2p+9b1S9u5cjDMIgxPcnD2oMaHkXQHLT02A2
CHqPS1/S26/vv0PBG2stMHGHlQzaSmBhwD1+gdyZQszDwHWKwM4i11WvKdFbR5DYr3eDmENxYu3R
P5st8RC12hAnqwnfTzRJPUHV4J3hTL1q3fBoeRNlx2NXioH4inu70qQSG/8SSB0Hbgdlgr/+EZQZ
2VLJW1kY7SEeTDxYxnpfpy/pHz4WUzYg1EA0xwoE1JNC4Nqdo8wfz7YXviH0AjulGSJ8ghAW9IoL
wCmT+h7tfddS9r6aSoptYGapH1UGCnfGgMc8YU4xBx40Atq32CpCqKYr8tH3saFJ/CJGCZm+eMHQ
2+pXO5e37exgZOUZz2X1dbMBvE3ZlHU8JK9h90hMkD4mU7HJvZzsjU8WTVOT+VnTGWeQBeMwayD+
jUqqtDDQM/x4QMmsO1XpdrLpR3tGCNQuTwtVAz1kfqYhGj0VadxwJPOjWskMCOaxOrXFvVIjnoPb
EUN2LGysZzB34Pt3Kr1qYAZyp13pPvW9ud6UxfgeL5fQzKGROxYnBvR+94LDqDBw5nTW28li1IpT
UEBaYJflBKBLlNVqI/THFpWhgcIOW7c1qVpy5rcB5uSkMdvoWgWjcXbBakbdiXxZRTRr2SnytGtx
WLppcEoWctEbVmA4IcmiYpx/rNv2LGxzZOmZntGb9uFV48Tu4pvC2Un/Xn8ZlcEo/JP1Xa4eUKDj
zNRkQ4hsSWD+X7kKs3JeR52CJyAG727BXLA5kIAH+t0W/STsdd2ZhwyoaOuCU3fF+TGxANgeIVir
1meyJrX/q9cdqFm4GeCZ3Fw6vyOfWeGEjfVsd8i2chfyy9UmTtvb04cvG6MgwZ1yxuwW/okSDbqL
QuHqcS2q2+fRYXZSZlLvWBKVSmBzJe0+/MNDG8upzb7xQq5KIx8WS9JqGhAUsICVTQWcrkLOrhTR
YW1SksDFnGX8utrHrYGjOJ9FKtIt9ZvF5H8PSxBIt/GMkbPAwiS6k4bIBUG+AA0PIwCBGuYOhyMu
ufoB7LYjKEkL5IswHu3xDJ7XG/E52TslpnzBB1gvT3yjhthNs3/cYC/Z2234877pisQP2yplgNL4
67iuIMMZaXzj7cwu/HBSTpVWOSNPWvejc2LI3AAK8KhLzlgGiNEpxgfCts88sBTLD7lLOizcV86b
TvugXNh5hirs79mwn6jrddrv7Gta/+5mC3tQn0h5nLuCeKpd+gg4bfHU+FSmomsmmSG1qyeGzYgi
VnydoKRLEeopTWHfimTLun6SsSJvFeA3AGl+c0mIfPzotNhkkumzxDU9XEmoIyPN1mOAENQzS5iG
TPlh+rUPmC01eFkxfTqX3K891GCA3t0m48arciZKTntZKx+F1Pw3D8EAJBcjwqwteQdwufzbuaqR
m/YRV73pTdypAqi8vXg9u2OkYUdbiRXPEq5VvpFaLgODonMDCORlaxni1D4ldYu9EXonKbemEHx3
nsmjjXG3psVZU1Jr/RmO2eBM/oBnVHyyhWXuVJVfeOiwuc06GluJ4LGRcs08lS+AzSin8ZHNxNZd
PIJ76zEnkDw8QpxI91oqTEoEzzx0IwzYWdwiJdsmBCSnZUmFjltWhEcDpKKz/kgbrubHQGjQUZt5
v1QOLFaCOg7J+WhrcykksvATTZxc3jA8f91SC9tzELcrwAE+PTXragdQOB/f0Fgs91YPx8PNySl8
alFVoz8CySyBQcRF3+9Aix1f+Bn9MIFAx/rCT1gu8nXVsW1O6CbJutE2Lu1HjjpN4tzHeJMxcAZm
0EYmIxyOu3YwZO85i+c0okO96wRhrgMVCD7KWn+g5hRG/iMonmSEX+sy1wN6URbNiE9mTyDAVDB0
oKHlzgsZfXyX0V8uAa6F5Tsp82so4eeF7ok9RoRWnJtlCC8rR8u6U6zq4vI4a+msuhmub68Nr9fD
dOsB3CLCxNlgXi0S83o0zQYQIJK9IYCyvsA3HEHw/2p8jrUXz4h5sAq2VXTTKXhfPGaN2obvZsAF
HA2wbmXkobDvOx1+MLNdvFYxi7mgasj9iv/AYKqGDvWFLQtgpD7RB4zQNj44omugtkN91Q1LShwi
exv+SRDXsux6LKnvnK6H4TUmMkRCWfPJbxDm8uTT+hi0iOQyOwiFrjDZw6LMHWP0enBq9jMGCbMf
U0QoIc1sWGP6lkSJCOdF/tLHUEsd8aRowaIfgJO0xpCMV16QdGA8BYUWIztfrHzIWt2VIvDHJO/9
vkskHolWGvpvIIoBRflRMpC/3PEpkDWSzUCSwjr5zHbIh6Q79WqFuykPKJsJ/zk++PiHkZr1WnEI
PafLHv9qxblRy+5EQRUdBJMTAPO4PM2AJA5wvXxprfra+6l0Dc06yIrDADuhJPLCutHmjRwqIwjI
SK6HWq+lGj1XysLydzztfIaJdjQtzkCj9S3khWVzD46LXAYkLsGRMS/pEdNtdC1hMf54LBiMpnZR
v5bZ69Or3dCoRSM9vw2rKfKhRqwbLYYg9uyXKbTS1s1TrTjyzQrRzDRfcWHZn08qpEH6saGhY6CY
Yj9bJNkuiYeb/w3v6e8TWUzJ9HuRPrqe3Md1iCSn3UBE0yf2QgZykC+sKzfzSqXxkQfvctgpUkvz
QU8b02ton+tkvZx9JSglfOA3qvC1kF2Q5PiFj1KJFQ+UuTo5njI9LRhDXkX+aA1gYvi59mZUfeKM
8xqqmTkDapwjay9QPnoDBJ5di1xc1UAH5uvPlDf+JGGaeBjaIHzkn5CI5eVaEJIV9/VQKSiRsO72
rPWuyZ4TWczPZztqFJJU9Ajn5FKzbToO3P+gwBU86qv6Ump9kd5FXlIZ9MFN0wU7UOboJZ47zjII
baAQkEefl+pVSJDVN2Cvc1Z2NVuhyZEJIFFx1RKcT0yZpqT9Y1mjMJLnMlGfjtA2OHXTldVBLHT4
gU2jXAU1NrtZjpuny2eop9woCZ1V04FEaVaoAMlJJhpD8aCS7pOncN26irVx8Ge5BkvS2VsNreUG
bPDIGUOWOyc7mBJuJlgNGixtNx0eDWU7CxCxVBRwhWu3DEy+NBSjNdY82cr26myssKp1XquEK1kY
nzrJ64d8hMdMT7FOlYRQdueKa50nd2yPeiNoUUo1m3JMdydfGHk5/iwRcBpkOWWS+G9FfVlKECN6
p9IpX65EnqIXNHGFLLb43dWSWC586cu15uJAFKKdDv5XGqQfYVnTeRmVoD/qdscZZ+0OinsbKejY
4kiJWte6BmNl0Rr4aL1f2AmnSMf0NOXhteuGQR+zJML6Bp5sFMUuUc46bsrGmtKpO/M8mH8N927q
VBQyzwMUCtcyRt7JP+UYpeRvm3AJ54uyxUk/BGnTeQX5Wt0Qrit5IiwRox8+lfQn5OibweodQ6bU
yVvCqBzhvk4YZBgNsCW46kxeY9bOQwq7/osWxlmAhMYlgMkTxwYjwSxSOA8q5tIaLrJxkQ3yVLmF
TJpgGY89rsc0MialK30jtjdzkD6bUOMxzKpicj3fBrXGZ15PwcuahRwqJIhAkdcY7GsREDS3KP8K
LnaJrThLQkp3qIIjncPSXw1Uxu7dRff9bnnPczNcs2VkUOjiY3O4RgyXf+BkXb7H19JB3hduTRAj
zvBK1aydbXSjmbgS5NW6UqqC1dJfVCWPAXVkPzdzA6o4nNCYvuxBZdbKrAuNBNbMl8KWn51aRfIm
bAi5mE5xizEwgevXYxzNOmrBPKdcVe2qw6niWbf1Rz0khITXhaYlhPVvkqu+wl8ee2cAg+vLhWgW
gzBGCr95Wn2VsgnfFReg19hk5AxCyydNfcPCeY7omxzjdz7BaaBsk4aCVyWE4YPqHzr2TS4BGsVf
SgHBb8ENRBV2Vlh19Jf6FdUlvTNYaajUeGx7ORqB+wf8TpP4aAPfmTXy2kRJvfZjLm0OarEOC2Lf
wqFNctyBpI46EzJCyAt4npjajVBF1rdj9RlfE5ssPV0PId9hJ5ybBy9x6IDUjzpj/cJdoutAWciN
UF3kRZSYuNGZs6G13gF8prvhAVasOlKdQ3DGmuQXypyNeMM3Yxe7HWdD682ueC7i3kRax0LTvdzd
s1MAdx0r2708fFJDDsQJOx1P+lauGTbaA7pBYRxeuPx7gjtFmuEjGNb+OxW27rhYOhQnVjXPGjgO
QgsJWizNIvEnbNJQi60imQ1V/+fVFAUqve26WN0pqyb1VMj3ILFl3LrnoWxYtghCkEJ9AZByiqpD
J66QqDux3bMhDGJO4YDqP/dECbdweAo1k9//SBpZdijgrqV88gwh5/Tq/uWMmqjQg35vnYe+ZZ7f
oGQjdvzzY7clC4Ng+rgEbfQHnw8dbuDo7x9/gdpHcNvorvq0TyYY4+crTVAB16TVGYjSD7SJJcFd
UcnYoxihSEZ38a62qDXSvchBoVIfN+m1EkWYYSXHJ6exCefXu4WLSBJ84eS+56jtzfVD+My4UEob
wdVU+kFZdA0TPO+uPbekW39CeU1iXNgNN0nwhggF7DygDht0Nbif+n2QCzaswP0jjy9cZFg09/aB
bpAlivMV/Dsu4ax+sACYpxNzwWZKUVKPDYJvp3BqPLLhudmw4h/fFx3WreEKjq3ZdlxMYSMUUtT2
afVHVWTjrmJ4p9nWwCZtP7JpOuh8nASBmOEXQ5PX9psyKtOWK3YpSKZiCJk+/RvwqtWq4tT/l6Gk
Yrsf8XH4Ei7rkGfHdc3MwOlEBG/W2zBEfxueXu9im1NE1EiW12b1AOdv3CX4+rvjpx25EALPeb/x
TVMjmXaXXf+48rZG4r5HpjP8wkxOHqCtDJveJ1kHG1ERTtOIzn2sEKowKXbtPCv3jj/Z6F8f70vM
Z0+z7meRcKxgFOuD6aSi7DWNQ9wESK2nfexvrjIYE7YevN6zU22KCfQUBfEjOq3fC+VJ2gYGqvpv
Tx2ooeU5YtKfKHwjfDbjNOE22/68jPUBfZ5taMBCcmc6lWh39OAMg8UJurDGAF1bg1XCMqTwZex0
Dk+PI6O/ARDyjOvEwX3qWm3oQmLL1dkDwJtca3AEQICthPDYKTXw0TTTMZrw7TxalQyAF0sCjpyc
TGqJkBs7cb0/ySAPZwNe3NIn9o12ScS6loXye2HYRpCx8aodIw5GuS2xF7VpMj9DyLqDFz8KVEkT
atvb3slKSd56hJKbDTRvGe+GZXd7i/V5hBuzv0JStiVXYuhix6cHgVB4c6q1rVAXcqFJ/U4SAFNz
z9GgVt5Hf7DDHdYMIiKRp5Z3EL1DyC47GSMYwTED8+kBGGcdAyq2UPiXsLlY8IGQxtfvP+hSomx/
aT2E4JdP5ZSzyr1MyrrgKjKdpOKzcm5G3qM2eH7tX0GGfSlDZe3ZHdiqYTXKG5HjRVYvAKGdu7Yi
IxdGnM19hx7zZB1GRvNcFLf6kJ6sBrJgoonXo0Ib5sztn+AfYzsN8jOy1W/vHGkco5ku01QYV67j
tA6FMSYD3OkAEIE/uRog156QG/WpB8AfImoV59oCdtsKCs45r2SAP24S4CMCZg+FxVQfvYi/vZqk
6oCuZbBMMElY12c965dLmcIvg1dvsR1wOTMLblYvohxAxNGodB5syQmcQKZ8kphgViiuAx5FcIVA
+Uy7506nNQbQ8JEYxNGTChPh8Y+AWV0htAke3InVK7AOQkWly5rwlCS9QLJxfAMSbn+nm5aMJ3Js
utAtjc/yk8HXUFDTSzgynzbK++60H8Up2oYVD9UF0cvMBg2mi6pvtCdQIuc0pvHKD55HwaVuusjF
KAUjIXZWt6J0ILxHdEoPkZE8QroVrQQgzjFV7aUu7RhkZOa7ewcjxSpaPUT3leyWcEE60he5AQhw
rPyH+Oe61Ee5FfLwXQeNe0TvGjx0l7Ii434OLpzzDLEzbtR6Z9/pM3q0xV1VLtx9RFV3YiMe/4q5
YajYx/yLSkBerxisDQuN5d8yhs755HA27TNW+wUetKEvStYkWmhPpfUDbcFF7S9nDRMLiYjx900s
xP9raStlB7lGdKWHsN3jO32wXs/VHg/6SQv9ffFC2tFZAp7Di7TZLZfFKsNCtdaaFOhDO1Y3bReD
bF63UbYN8qaBSRUvvlWz2BsA+yhTfm4bG9prvbbxxZXnVKDwhgEFiiejxeKbbhinKomYKtWTXu6a
E/IMi0Fea9SaiPJUDd77WK9mU0sVBLYB5i3kgmCqLRKWQdGc8rh/ZFBzfPAFDxAD1PNf0DpVhy6j
4d2K/iQhw92uZD1dV3ps3tVFe3CgBJ/Cm0GQ6bo4EMEDiDcsTD+ZU+Q3zcnzUwaPa9zzw5t+MLh8
ksyFwAAH7xFL+5jB2jzZ1c8YHKk4/YPOOY4ufddN0mXI2BiAtS4YrUeoJ2tz6MJ4hyt5WhN8XITQ
UPGSK04Q5d9NIst97nG30Yd0zq4AOve/BeqPH6eudh4bV8OqX0sB/3Iv/0+X4+n4HDd5wAu2ExP0
E3n7kg4vFnn37k+3dRCSf/WIzvUEz3FL6Jp2DjuE2PYgqP8FtsMbSX2JiDmOf0KXmCSMZx3sgQR1
KCmUcCgJC7Ay6M5mkWPT65dIOBNYWsekAkhWTsn5GijhUl/DALbDUyownQYAnctJ64CiuJodM8jw
u8OOHruRW7RGtKdgils5NyLtqg28mBWGxqc7qRvb44xzzZv74ZYzfVLwgTPWHDQHjlHX42PJKogz
4ILwmwiDXTlVIpLVmNjPg0CuSEavEluC1MMiM9uhRo1QwiWnNgR47u+tczxbCAisSNgxxo8thSFC
frJaH6TwQpq9Zzno8HrmqwSqQ7vpE2dicn4hsp3G+LSpgyy90TuJ7P9CeGplpjQiK1k9NIne9THU
Rt7DkiwgaHxv+kRpqeBTm9OfaVNheawq1o5ZZfNAdV+YwG8cA/4w0S0TTllyh6D4yY1MMtyG1vXe
qHG07nPy2oeWxfcRiKnbwAhFTuvjfZeaXbxe2Cpd0iXN9SzLE1ftGuLHZ1nIA4/q9QYmTjHaWc71
72JW1LY/0Au6T4ivadVAanT1PpvEXF53fcI3+f+cvjXyWDEjJbOZIPtilCjuglsTCCzYtHghfU6M
UDyn02+0169hyg8sZw1MsyIyWCB+EsQRvIdtYvwT2TGXr/WOUlmdYBcX26QZhncnX2JSMFt6L7u2
EoqMC6Le8B8bgNAjIEtm0eeA1hhygmViCIVX5ca8Ql2JEmUw9ytlTbHs9ob/ssqFENuLrmMotgxN
JfRYf/MYQD99eHrXO6QGaFAF9A3ejbtbmC7fD5Jaz0NPm5EtqiO9CSqJaN2HWmFpMtmHcFXwnG2z
UXVdLAsoZYQ1eTyYFBrow8sOb+fbThMHQP0Ur7YVZmbM1bqOQp7yguOlmfDEKDSE8PLiUtvzkmO/
2jVf7YhLdpOTs3o0oUFTCESe9/R8ienMGuApTlliq7t+YyXrzyeUx3aWTpFPyUfXKP3gfCMcs8UU
uW5Eru1pzzoCoRSremD9Iygos6hqTE3E3BSYZOaiLRgYwR78y0KFxEOdE/I3q43YspgGuPNU9Bi4
7pmxv+bRBJMr4LFDpuvvI4+EYqBTzHce8EXTUfOeqfpB8E4rhAedkfpda6elxdrVoFgPhuKbyDxG
PqG+5L6ppOlpdy544vPKgUJ9krAeDoTTIgDjhD9Ri/+uiGnsnKqmkDcN++StRIcIfnX+0zXVPaHh
kp/cpBe1w9jyyzV7EUslNPQ5AK+5xY1b08TTmQ5Am8eHuSDeK8cF/2Mkw0iyT4rB3dd53jwTcg3c
HX7SN07I/a+U4rW/OvfxC5OskI8bx2CRKspMczMbHpr61YDxCk87SVQ3xggD8cZE1+GivqDVq7BQ
Iv/wUiuZXN+zj+dbwiZrciJ3Q88aU6PnFqyL+nN189kuYAygm1XANxVH+3SefP7E/mxfd0Y+m+ZB
nOxUJSPEri9Jc6ZpM+Uw/qiSSMetQ3VNEaXwKYA/0SYNxtDIl6gWvIl8+kJbLfZ7t8h6EfKJX5qh
6ohhx++hsoEJ4sTDhFlbi9Z20KaazYsiTmWMtwGPmz4LJTrKpW6qvHLGoCanuCu7w4S1+8TGS2CG
Z4AsMqjVRoW40o/26qs0OqPaB6KZBQgIVAXVtv24x9wXpBgUj2TXchcdObNTaFvh5qeOfHtagT+3
TWA7pfXor2WEqQeqpmFZbVA0GpsdxprCp3qrxfpZ5Bzhx927krIt9XyOSSRGQep3xpde7QvQTdAO
20NEXUR0jVnycRDqcwEygrscplZtaOTZAbgrMmeEmJcTr4x57czWHg9+43seUyXdllwL5wQIqTYH
SeuNEgPEVVjQzujhhnXjFadImXCVuIyuB/9czuPPpsS1Svjd7l4H3YOf/RQdln2CnpFYTbt6/aVW
FjTF31el2/UcbVtgDD4vG8TIrKaSuAjbvpPpgVVbRp2pie+LWHOTczH+MVbQpHlp+d2SdxR45Bfw
XBmR+WusNf7oTOvmoPSjiC/XRaNzTpU0OcHDfj7Xt56ppxcZ2xrh/EQdzIFy1TVOUn0GPJ08oLE5
Yql+zq38URd1jWpiPwpWW7GuIo4Cv/IFLJ2x4c4IflSA6ZYWC5g7Mp9N7J+I1i8SvfDlF7J0tWZY
uPEezQFns8PHy06X36aOEUQdK8PeJs/P+10Oo93bKw/DjMvnrQ9BpKX0PAbnMfNo0AoMb6QMO2pR
eBlkRCrmXlgbjfNUBr+hsj4dUk6m7PFHVGkIA8w4Ub3y5UwZwEq+Ubw5bAwjX7FWf7dJtzDWa3yN
dtHMEDrNJ22uceobCeQ11UjhDdL5jwC7xtwA2CMQ1JfCY8L4e+eTs5p0roarwsOnb9Edme8qKmtb
tEb1m7QxOjJ5BELCzkAUKxmKHWNJSeM7ACzHvdlNQPDebIZtBSwzvDq0KBley/FAlOo1WEjiaRbe
/JRNtEHoBiNXPoWiUObu9jRRWedrrO02PkK2Ww1iWhh8FSmKv+ZEy/hmiZZURo5oDOCkZuZ0aDyx
EIpuEn0Mksm2bPtjJhcKe3iS74oz1BJy+w1vthCN93NXEl6Vs1hC0dQ/kDuefzvol25wS9ouFv/O
FT6Tp2/tTU6IxQyPfRIcGsg14UjktT58uNk/KvyNERbevqUVDDYvg79dHg+lzZ4XPLZU7rpgQlhz
sIbJi4aCWF0LFgWckOdkW7Kgdu/BruNmQwcapB8dnn/wck25M82u5cquXc2PNgG8RyTecIuE4Rur
TL/IfhecT5JiqKbPXqulgp40QQW02vQym577QyGVi4tfboAh16PyIXiycdOc0daeQp0RbE9UmDN9
shtg++tjG7lA4E9fBgulxQYZdh0OjZDwJEgqLoQmDovHlPSgRbdPtGrtusANHWNN5pOLnnYwwM/0
AU2YPXgHl2KGfaZEHXmJ1ZVC3loFAdFCmgUaxBtPdM+TVvEXH3yU9QbVXCRCmgNhqs5RvlnChVL4
Tl0ir2WLml9QAC1tCnDr8tD9R8TjPC6NRRvd7oo0xwyZumG9QX7fV7RG/hayXat+spykDeeMGr4W
pryJkBJX2hr1HKQa5dSmmsSmrK1kRITrMvcZ8QADO9ygxTn4z7FUDlxBS41CpQcwrwLkQI/wMz6e
5ht3mMkI5yOumpgBTX8qn0pqEBHYULl99MPsW5VYCPyKfZ+qrZu8ZjtK/QkklUipVVTR9AmoQ4Bb
SLYGypCC4eaVV4BrJPsYgb5wx+KwxLKhv2XHxoh51i9YpKnRSV4hMPi7Cq/86yCEqWj5ZNQTGEin
W5WRac8bFb83mXs1zCUlSK6Ho/hsG3GpTvPuhPBLYDXVpmTApMPGrFlEDV5Vu/wsgLvNxkFjlko/
NV/KKctVAwfH+L9A1Z8yKmZMdMuTwh8g2V7eEkQEy+aBalAnNzSfW3ylDwBGXzUGH7V3EduwbPnC
x1nTwyUYey1rGGlfe1kB61xkBl1FjMAgJ7kZU483nVJ3z5EIMlOHTNXLLMWYgO01W1mts2uzW/T3
pmdqLVF2w65a4/f1tzX+oI0qmQDu5XlEen626ZdEWLobJCFw9eqpYU9Y12R8EUu+3Mn6gIwGFXHd
CD1XVb6p9nIVtMfxG3vaP5kO2DE+KlAVKttdZhMQhNzVTM0zRFfP/JUmuaKgb4UecnvIXVgxNIZ2
heMlnYSRHLUDE+ftg/UHFnAWISeQyEJ53BIa/Alj8MljJcmSQZJU0PoTxupaad4hpc9UHaLU5ni7
isSCDLobP44y+MxwZNetXMQK8U0WMyQBOz3sCVXQteD018zyBfH/0SH1zbXmVuRlhbs0y64pgdXi
4YlwlvHVfBMiLClq1qh/Qr7r516Z5Nwb6O+/oX73DJ9tljgKIfLCnA8s+jUqUAzJCLxqG5VccPee
PA6wPTCsVCGX1BPYtcvy4fXVTAmhJW51ZQuA9A11GJUz5d6vsYto5iDIcKHUl7xhHivFeQLMsVV0
1X9V4TVWfmyS0aDKpk6xlY6icTB3/pIe61Sw5SB8wExSSzOuY2pEcXVLyW8B2UzstteiiT9UoCcs
0lxq1/FGxj+LUlhqdnhJj5lNskPInFuz1Fi7TKrik/HozWVwfSCFRUgjWANChX7EUQkn0AAYInfc
tma1f8bn+fpY9nDs1CFG0jXxdDBmPGz2SkSuJ09Z20YCrQPcpTS9TSjp4l3+Mnwx5Zf7/uMop59M
mR5HX+5RY1HriRK/Yt0+5/2y22/N1BebgGKicH+WtS0dj9q/mnPFrEhK2e7AHhvTplON0BIrpL0V
ocaZ9gGvg/VjABXV6rqQRSpOCucPz6L/nA9l1weHPgapZkEMNGLbEVr7VuJG4QKT3Pm9b4qqygJU
me5SAA4vCzo2WXQcix0YL+rHhfmE0osX5oxEalSaE+idIY5pve+cs+Vhhqf+kgnnYVevmRER/f7j
ImicRqs4Gj1sRH2vkFhopuEq2ew0O97zxjmMQMmG8cJSxQps5dMQhDhhfPs41G/OUBM92V9F7NMG
QgioscRF3vPUgRz01CfO5pKb97bPx/kKNTJyeVyHN5tjtkaHm5B7htD+rgvt5O7qjoN7QndduDGR
yxf/QHSa0k6ifCIdqvZZWGpooIzfJoaPjAmn4OpFfEoMNwiRcpDkKz8P9bSFytrldpveeBHVRHns
v7jO2bG7lG142Nm72pTkjYjbPAVkDmX46hiCgg3RjLXh+TR7R/R+FOcRi3R89Doe3fx9aPgz8ZsJ
MSkrIHP14nqXlnuK4OLcPcboJz74wuCL3zghuWixGuyYtZKNRqfr3GK1kVUJePdGpmjSINa02pKG
xZg205gsXu0xrAKuHmLtSIdF3QPRw0Vk1+fgrN5WwPAZrgavDFVXTbDi+j2czyJBzPwtVKYieoWY
wNjo/pex4kefYBb0YMm2A9f8XPcanNFzwPW6G7PhYSRvCUC8A+bQLE9Upm32xd7/j5x2nNREcUZM
2UiH8O2CmJ0dePYDIY1wn12Y66vHKvhfOPfFedrSOBMgSQxr1e1M0gPWLdHtFSmM1fUCAov8/weW
1jH8wb0KzXBCdUnQhQHhdSwzVCXLg6d1e2NRrjEx/j1IpvKz+FecfoR94rxSA/tBWKTdm1mZzp6T
cWQde36Wjc15dI7Or7ayc15NU00vO27lWkOQz9t5XK15nybcYSfYRH0szt33jhU0qXj49j7L4/uG
pez6GJspvsEecpLP/LTYfJBMEUYKZxyUlIqBEZfaLeoDNgX8GPoJsTyKIsvNzXKeU61YP732Y3tK
4+zigJgnScAAV2vnllTEaJnyFV6C4kaBtiRpCO7cE/8nknTbejPbyQEVskw3KQAL+O4yhFk86NQt
O6K659TI5ApkgQlJiB/EPv7WyL+urJxrNgqYyYT78Ex8YZL+LnHsDOdcmoULYSW881O+bhYrtFOK
o4dptzsirDk67vPlUfGWfXgWMvKE8ZU+KOLD0lDXa35QzXNMyDo45W7hJbIvAvir/fetIaDojEZi
48pL7umTDTwhhNkH9WGQbP1O1+zIrFr+L5mTRICQY4rbIB/hAkN262cdrPJg/tRyuMid33fQBAMJ
3OpiTR/5Su2ZlcHMCm4/s81ZFQwBrOVlqQeP8N2mP3bNigVoQXLdt1+d26NZlHPnUExYhovAE1go
YfRVomBMQUTZgv7k12UNCBKvo+W9zmbcJiyjpqGnmFiFIrHDhAMpCr3CHKqDFHDd2961kiZjhwiv
0fzElWB+FZzL0O6/MAAgdX/lmQSaEA5ZMkPd9L+tHGukULJzMj62DDqYqYhOORaIymdpyVxnlxCC
SYLtJO4hc33471RxD27p0VRDUzh/qT/3STUY1RoAYD8Gwx+6tFvRzQ7berj94gviBwnLgAcEhlm1
G+h3/ytj3p5zv9R3pNW6R228mPESB6SgZGJTWzAz0hG+W78y9KOj4H+qvVgc67nThP+lrpiYZPrd
6Los9Siu2WL6mHEk3GvDlwxPtIGV3mMTCexLG0vOx6zvpmuYMWsRuXwBzfiEfo1yGPN5TZRdSsfQ
VsgaZshvLqmP7fgEIndJPbq0ceWJBGkj4yZfv3UdXf98SzY5OHudS01+/4d5X0DUYjn88XS4P1fo
lB1/QJfdaPBoSW3zYTuSZoxm5mjVOjPesodm3aXgzY7nIUfj7+K5BOmzfMmMf5nGGry6sbvst2Ot
lfkbiQyxxspc2gW78yGfD+nVwWjJVZgIoGpD2wW9hUy/pTZvu9d4buOvhilWPcLRBWTbQZAX24yN
62liQx08JgfPK8mjOZ7JVx0QLudJxqai1VLpk1eGwKTtbB+K2CZp2J1NlTXQ47h5PD2MvYoaW7/h
uP1R8Muu7hsjkXNDuwJAf2ufWrhzmGAPQ07SPZwd38LK4NEyG8cJI8vngpvTmp37UKWo6vfHBheI
puqunL27uchAFo6KdjZXU0Mj8yEls60qY3gyNN8nS+OtbEkgtyH4w9UAw6/csUhLH61EMIpIk+m0
O9Ysx0RDuJb5DJni8hBH6C1W2bMKyvZfnfvfCP7I/Zuq7N0tq7LISeyQgxtw2zOkbKxsCg+GQi/f
D8/5oJasNF8JbcLo2JIKhgLpudQ3BdYqnaw1tuHafY6xl2lFYaMb7y6VowXIfkCr6o9sw0DBgICZ
C+voE5LANLN1XK51zbDw8NU6yEU+yNBZsjpwd/q6g6ihEkHgMwy1XGaZ5rghQuuMmfF9a3Ha7uDh
8wL+HYbSjd1YYb8bjvyEug26qB7drJIIBJwGSboHxQkApQ0untofRIGZi0UAqNuYs9Vyt9+U1JGZ
ziJ60oSSAN99RxnzsFpYUBPjTr2osMac1Y8VO3HgDGWtDWugvokU2RUu0GWkFp8yP1poIIodD2i5
pDVWrcNl6yCUfx623X+aIiEl5SFDQIS3FfkP6WT0V1LL9YxQ/VZsr606HortQUmPNu0h9oyrklGW
43v9vqu3/UT/yODz+NXzs++dHKbtldMmrgnamQXsalDZT3guVcvrUg0f5J8LpqHOax6Z1ribtXGY
vtnvOwSXdrL8W8p0csOolEEVV+F0qK6wH/Iv5nU/xh9x5CMK9mJQ7YCpPfbbA5AfINQuysHh9cpY
R7Y0RddlyF7zyz0MRuB9hDG3ewOjhxrxS2kji8ET0vMZT8hAiX5ci+ha0n1AdmPPGHZji33qoG/+
MVPk0pYVUae9K8mbmur9A4iL9PhWcnr7oIHJ6Vc6esKZp0fpa/qPTtYCQkHTyShXy2XRSJS4Lnwz
F0Vol1xRtXDiWUN6/PL9NtLQtzh7IzmLE9KtkGPF4uhxVTBx7uAbdbEdx2pSmJnt0ja1Km4HP9tj
eUVMTRDkMs87PJexNMFmGJd6nm/h6+v5bXH58Wj3G0aqK3cTMLo9Jjvo3zaoKfpZ7xOWC1OApxtN
VLwl7HG4XzFjQwWEDv9G98VtHNulVlr9yfCg++REuJmQRH5JHRw6Iu4ESz973bcgjlk+XGROrg32
aat1YbSc8B+Z/QqfW6o75KRPwl9ILpvwDADERASRh4dRSUgyKYi2AgXqfWoyWN8zhVO3JySf0WeL
oj1PvUWL/2yO3+Pzb0x6M/BWbD4q3TUOOi/m09wbgfgAD0dT/XfTlgp9yyUWHbqf6xxfnZXH1v6v
/xpmLsyL6v9UO4fS7C+2kmbeWgg08907O/ezXuI9x8ZEEgoRFY7GjAFcd3Tuk1ErAGr1jBOf/+b9
QGaArCxxSinqu57bYLonTeC6Viu3YERPSr16sv+1v7yvh4k/lW9kwBXgnOyIFIcpa3qA4RRGbgzx
L3nt5Y2+4lLc600yXc8G6JvmJf9oXFDJQCUzcokEV1WGYx3Tb4sJ8rVhSIeECKVWOxqxUWkinfn1
SRXH1UW2kyxst9+MVctcokwJY1awXJuY9NE/HbAAZviMRgBRnRwTT3kOTD/sMXHxFp1lMF4qNbEF
P1j3HBoBnEeaM6mu4yp7Z1es6u2Neizp7OT6dvjkH71InXTB1PuJY0Bjw+uj6bNSCBjJyF5p+c2k
gJgnZxOMK6ZPcV1lFBwRBVQzEJ64jAkwBf8dl+/+qXVN55/cMKmkJeac0TxdLF4+H9NFfUzwpVXu
gGn8SyZCn/XdHgNX3p8FZqevpi2H2Pnwqz7RSdSCmliExeBLZ0iz4YFr3/pIDqb20c/Iuk3wu0Wg
zYOZ/VoYcPesQtJ1/5OHTXNx7qwh8FFgJIRM2q0ZoGA59w22ZlTnhB7AO42RzgpPIbwd2etzUC6m
yHaG17HKnHY4dNV0Qafz/H71lsL+Z9gHoZ2CNi56UjtQG9PjoR/eXNMbRLy/RpL1i+5dULgNs5SK
74HoJdKjdTkqeM6lejZlnqcqel6J/nODMV2psk1beVFIsN2vHJF3zSWLGCP1eRQz3iAzNidVM+04
pVdPqeAXA1l3doYqIi53v9JYYKejChjZ/KSW2XzYWTbrBITVPsDC8y5dY8rlQPS1vdO7TjPdf3ew
Wy6Kk9UX9sFgX4Zlq8ReVcz2lQ8wzBm4XRFRLnK7+yU+cAscalrDHDMeRmV0YueRGTYZf/Gqnlp3
9eRcwSGIrOEYz3n2/jtfWjEtDhbQD1c1Sw8nlm++1Ec8Srk9TGvV4p/gq+c/ef0YeI2qpTtB1T2a
YlgZon0UKLNuCJysUQvKg3Dq+Ms7kk0FivZ1Uj4nqlRcs2heF5bkO0Bi4s1tCmX8eUbtC5EQfzb7
KW5gcl7qJXc2fNcLinXSzDGlMo+qJkYQM8qMbtmm/EGJ92+ArhM+4PfAUwEG5KGX4NBVT7ssmoxg
cd6kLehvBwdnIPBocDzmnY5xCyOguF1LjQA5g97odQA9ohsHMDxHtfDkw+NozSq393k4Axh31AeM
th1XnHRs3/46OZh2oviorgq6wlEAP+1GxfYCroOvVm0bhUGjj+RTIwqkPRU5tiWfu+cYut0OUAe4
LnuAB/y0eRlxC3QwsIZTFcnSrdu8FSBRFK6CistD7wC6ISPuGr78iqLdMhED17Fr6oJwW7HdcJQC
ZYBh+gGPTKnu27AIGOTPOQBUbPoKBNR7gTn6ULL1J22QLuWSGEGwpY54TU3o6MtY4dJ+xVXgrJkI
CdK0NIHriJfk8qfoJFnm8FYPEDTLH8HY/6bh8e23WWqlvk/fO8Yu0HPVNEYL9dfGbAa/quvyUAgC
GZ3B9MomttQ4PMoxDq89K+OxwA3PB/GhulkIIFeG5M489owQefC1vsPcvffy7wLNb3EYjoB8StCl
RQeW7BFiDjst+ARULx5Ghh0feBm3hhp2asQugQKgkELtXbG6IAdtOO5n4CVoZML6yUMiLkhbtv9V
7SSCfCnFgTaKuMgYOZcCI4RiWWgKdn3OdvHmQz/NTilJhSa5djUXBgfIORj8RVVrZ3nWbJbRPc5Z
Z+BzLoSEwLLbc+w7bRXUdjskghd6DL3kyE+U5zmwF41/vmqfg0JxUoPQjRZAN/R1iql7Zt1MylBE
aT2l3yffKtqbN8JkZjrpRHHT44gRLVq5wuIhzD0jFzbF8U+vk1gajN645BHbGwJ8vD89yeTtO4ox
ubab0Q8FX0Yj+MeByxs1drFC6ftEm8EOrtVh1zrLvzt+ML9PfR5ODvTVlMqRgdbZLr+XBGFNuV5J
T/A9m8c5Jpn/G7buJOuTG6v5n7JzG+2JhdB+Ia5U0nOUdScrZV2Xu10aYkRdgJW616y14Q6ZTFl3
hY4hZN1uvmE+T4y6Zr7JudKe47wG5Nef/sOOXIdS2VNeVHvBSzC3NgeFl3NKLVJMLeqA18okTva2
Ne69SCGx3nUb2wNGQfJEoiu4uIQ0gGLHprKOMM6xQNL5oBijCETx9k8WrqiQIZ8Glex9Jvcv1YlV
7wU3TPD//Qwfee0eN4AdH640G3jBrRS09RmSdpKIJz8XtJOuh0tIOPfgpHEJF6RFdi5LERqaruVL
2vnwxQYqGrTSsTkBFpX9m6c0nl6WSmTe1HHqCnkEnA8bpfCL7sK897UkdP1oelw5pOoKSpzI9ArT
XCZxZmLXfx9t4ZSjjcGWAr8VRGFekKeNvhwIpKhRtxMUdF7iLzWl8GEhWzkLoVBoHs5+E8ZgEG/T
DKDByHZe4g5MJn28dmWBzeROP0BjaYbwi1YP4oIwQEUGnDnQn21CaPhCXMbA6VdPlxiCI6o1ADfR
/49qIjoMR4cOsV/2xIjit5+UePtH0Cj7u9j7qVksn62hPGBUyQ32kt9g/ZhtHcm8X2F6mBqfL2ZW
QzfPlqc946MbwAO+jkA3IVKQZfEIqddIHvmaHPyKVcfmiEmYBSOmJvZxUC46iMNcHtvQykreVkh3
UOlCuSKoh2c6WsV665N2HS5QtlwxlNmV8cXjy2URvzkOYBgi2G33UV0uZ6JqZQ9OpHAJHjChCT73
YOzy0VSXGF/9ZaBwaARIffux/BUbHadAutYQZd9lqxZuotmMO2EkyI4ckz9vbSiLN3PMLydmF4rq
BFybD7AR3k948d7KPv/7KLD6yCNwI+2XSoXDuMxpvD0T2tTcKSfEWgq4weCycxXLENO3IKYRABkF
aTnav1eq3uufapb3lJlEgpEVU5FYRnyd8gLFZaKVxziJ7kDqhSq/K2CFGkGuNnZsH7G5tt5zyhmd
kdPPHBEWh2xE4UnYGlB5kWTUdC+dVTljN3Y+A5fvP4rxYoPXeHU6fFczF1ucXviZPz3zsAD8iFBY
dvhmgtv/C8gGS6sapEOZBPii6RfvuudsH8JAOqLudObtIiK5XIThiH342SFrdc2WGKQn+4eckVjl
C6UaSf7vUjnmRIat0fzi6x6fDblj0N8vRbr550WMBeH+N8XakkTO06uITDF8eRIi1LLlNC/s4o/R
5qeVvQ6QEDb5G96Yyc0vp376vKZp+wvoBLQqc/meP6SLbO6BVed0+IPF7hDnHdT/Q7VABcLcQywr
zFhs71u93dRySixJGRRXR5yUTbJeqqC+XCmtxv9BZBcVkvZZ/TcNFnXBEG3UNukRQ5R/cARKh1Ru
WpLtsW+w+uDaiHIlvoqr3Pc26qhxEGB4UyLR5YSCM/IF9oJyJuTydk8lSMYEfGgqKVk2RFf0RV6P
rmxuBIqGyD86hj7mgAX8yF4mVTxpOCyP0qmCRk82vGaatDoZQe9cf9EzFZyyOo3QKqZGzdAAeKD4
IBNkn62dMXR498igg0HKnIVtdIOGEL8LlX7IFM/Ga5M5+Ewc9+xgk93DpvwvpK9PR7dKNHd3q+Tz
NOwbL/kzMcAHnjpKgVKO/Lza4lqn+qgR89dbk3V75FaVPhMN6WXHLXiFF+5IswhjOUiYjL8ycF2O
ajwpnRr7VmKYCwNO5d+zWuT2ylJEixY8CFphN/phXcvPx5d4nzBLOiBvnwKCJkuGf8aXbsAPiTgK
ZPH1IdrXt5BtI75JWqM9VHmXBwdN4YG8YJQvK2L7cgGysZVaCXjm4XQawoGtt9GHFEJ13ZYePeFk
8JzsYHis2UbEM2xG7ksIa3t3ucZ4g9v1QRzC0hoH5zv+2Ma1+4o5XxEmebck4nn5bnzRStANTkmZ
0KhdC8Kzy7cB9XBGMM5z6wwowMdU0FKFmfM4WmNP/05l/YadXrUqR3K0Z8ZDaQt71dv82CCTz+d5
4+/KGZtdQzRDs68CHFdrXkN2T3KgmE0+DlKvYq6b5FtrHEg4d1LTtP0L2jw9oyr/hAw3GxiFIlkd
7z8AiQRi723jHX1UeAPbkuUdCeLYz07c7hY2oEZ43gol8hldClAKHZ8IKvsFUhXKWDZ2R8uqZMoF
UX7Rezj+8w5Sw2o5IJjjkVCCKXVka3SxNvgMH7rtZGZ6o6jyTo2B+8eOtuONjkrjcEWclJQO0WU4
aBDLuwBm/W1A+pbzvMyTDpNm770Ovx18nNDFEGDwOMzf1jjmgkKhAvFoX04odxLWwHTBLREutigE
1xnidLSGqvnv/L9s4SkH0sLA03ThtI9DQzX0w52iCY7Su9nwYPfKoBrEqXmK0WAFHW5+hto7I3YH
sKiDv1L73A0XBrvmRZ0yf9vggGqeNLmiLF0S2aAKx3l2tChqakAp1/EAMJ+bM1exh3lUHcWpGfWU
9zA0I6vxB4i4DPGrk/FeWmMT3FzaiG66Gpqxc+DHBrqssPvUf7uHxpUIBNyw8FlzdgF7rSVjVh+X
1RRPqY9IqU6mWKWFaNdJxsn5wX/tLyLsbfUxwPXclZ/NzvCyutJLzeMtrSfxdslEx4WTc6WBswKH
/aYDYh3KZHHM0ACzEIacr3fmp5S0lqUfgVXQyO2XqY6gyk4wCXubA6uEk7Z9Y2z0MqoL2ZdFvUrb
Cn6w64QOhZ4gI4VPO0SUM1B4Pvq7VYpj1ciyzu7DA7LweHn4mjBUuJZLNLz8P2h2NAm9SxYY3pbD
osGdFdLFWSuU/Z2mLLhPGuRUg4TO2ulTO4KdwXdiQtR7Xq2D2QLS42MYeZRrUdgpuF7FK0b8JvxE
xs6VC6WJSQbLq+Ct+E911myy2947ZltQSvG/ryrSAbUztZE6imGbDFnFdPFZZHJhfQRoOUDol/41
uBECTZeJmf3p7JHFldVzYazKqe1Ljd2Hla7wAr/A+bkXD7Sol/6qhzw9+woXLY7ef8gbJkgiNFwg
Qsyh/GtO13N+u+UpXKWtHYw9DVKHMm0e/DvEaR6Ki6dBxMjfsq29RIiU8WUxO2doLXlxGnQTvQbZ
tPC2vSKqnnaqUQtXwrofr/9TTHeFAZ289VP8ySd9XBW3yWCAGIOSPdxnz/tfSAma4iAr9kNHPeZM
G+7517gwXkPAuBdJZS80JaHjSOV79tg28aQqpH1C6lsJuxmD7GT25JQRsxLALjnIFnALkvn0cu/M
Sa5u8bGXu1UR71DSQpJz7pAfsuuY9bbNx/WNnN+LE/jJbI8d1NLztxBly409QUJQiD5r4XUk9EMS
6k6b0j2mjNLlaVQMcnVg7wmYqkc8EmhOkBGsfY8iXZhRqZII4FYKcQqhubzNltPDPBGkTpCJYUlM
5QroZSb14II/ylRfAWZcF6q36sw6i4qliwFC+HQLhCd2COwSs+Yk/6KwA8zyctr1ECpE/sdOSdD+
u9xw1jhK3s68qdCYOO8H/PASR+Ee9c9LJYwNKCrXVPs3VW9cswVegYu+PMh0YpxEsHOGlngdwaAa
Zto5ERxgjYP+5NRVyDAM/Qq2ziXUEcI5X8vYNgmdeAu9AC+0i2CsPUTkyxprkXQz5IIiJe+W3m5B
aKyzIfu0+jhdUiOOKOx9pFzQIxLMscNxM/YtjmPzuaTkycypiuxk33iKsp5pSAA1lCjhGwoThiTL
NK1EZARsyKbOgVEoQfV11+ewU9rkN3DNStUHJSNijE0vzl7EO6dYQBVS+OnWOLtbPY0x0jAQt++q
QS8U1mVCe8+0H6szienLej5BO/67yty8XD9SvcvWEbZU8l8WHUBYMmLmXJrr0juotTZyLbjWMl2+
hLR5IqeTCRXxcgYfL6EqM38kHCtI5v+Ia7d5EucSFZdJ/Pgj9siVtxcko9D17q94Htylc1EkKcM+
SjFW57U67ocp7bYV5FybwcYquSGL5AkWui6AjH+PB9qrz3t22S6sAuQjjyq/tmnoRuqGZm6R6Siu
9QWcBzJrv5Qzf+jTVCuIcVIsYWatxRORtkLocLbkxhw90E6E+go1cQLrQtTrKVGa/wKYaP0g0YYQ
z0GiIPmEbFgTMILz+NqDG4knS8B/OgoHcxie4C8o8GSqXg4YooHdb03low0gTszVLH3gPN2U+//H
O6oFpfSBdFfSHDw6Qg8tefV0TxljdIeIIHO/EGnTvuCO/g70Mbzz3eM1lUzWJDKH1okLvbdYxjQg
7FsPJ1ZKxJH4i40MccuRVA18scUA04cMoOtwN32EY4dm8KVThUxkJK24Dx1YZJNpgkOLHXjASn9l
NZTfEtx7PJ50yeQpWWsK1MMQbpb+2UasghQ4T8XxP+fGBTN4zH6TMgjPSelxTm8B5I63eIThNW0Q
GOU/WgjjyCx6itjozP0SjLzNJhReukUtWcBOlRhe7itE6WzHLdq+6qOrKHq/17jhgkVwE24o38cB
s9QUvvIJi0Kw0KkrUlHCmewnSRrrQU1v2a+8OI9b+3OluVMavmMPmUM4HmVv6jyr6muX+XnAy9Wh
I6i+gBM6IMwW2z8kf6EE1cPlz7RId+N2n1bMDtR49OBppSxosdHm52HXzd0ahVDRYMiRaSIe5ohA
ZJ+LnNRtaV9orphK0tTGRBCFwG25PrIZRF8WPu0ZajriOEqsG0cBsUvZwbJy5B1mVFzozu1nshuo
MLRLISKrVLk4SICx660u0+z8oTD4qYADXbMNMKrz2O5S2Y5N/wID64O0sed626ZqeRLLuNutZ8RR
heIvROQMfb2OjctSdfGQVf67dTBOWLvc2hMaTys+eBgGcHQVwEabc6wVn73qQxDpDFxUnVH/QNL+
arff3DZNDYePosaNIKawfqS8TGQ1RgRBY57wkld6usNBurgw4qJAIOstexHXQBZRbt2whECKPMOU
JySUbHzzTdQy4MW+6h2AvfJw38YLmWyCw/xhWotIBJAChxHgkdkDUntHC4dXfpHfVkohIn0kGjnw
u9dZLj8OLEJJ/aXdIwXNSsHlz1X67XsekjhxlV8Qg+j5NkwIPn7ZfuwCMvOCePCqjjFkCjf6vhXx
D0hnI+euPbYxSiuR8uWylEgjlji45oO9/3EG3TmAUI7mNFj6ZVJeFqiQ5UrMrFKRTZXV+3IKjiF5
tBK4PmGRYgwLO4+YlmDs+A3JS9x1y8wgj5kxwO+25ROxNHVco22PnQ5P6j8bEt7E9Vux0S5pvZAU
gh9k9mgUBNEBjfZkDE4QTacZVz6IZB7FS5prGgZKdmOm64UrDkZWtZkEBdJY7Kjosp18foljmgz4
1p7QkfTs5qGfu7JO4M4/SucAoEVXD8y9lRolgjdmiaDUZghCO6Tjy2mf88maAYToV1heptYj0SZJ
ECgHDw4c9EInIrH6tnsDbDuuxdrs/euTy/I9ANd/wmT9NdG2IdY3R6dX6uNCJhQ5gjsYacNWWL52
Fq8Feib3dtEvj0s1p1BunqYHwyrfbksSjDp2CLicqkZJMLt1ZKGEMqfF4m2EltpGRfGBS5TX8D9U
n6ut05ovheQ99QnxkVoyOqQ6c8CFBEcYnJvbk4GKV74H/vEO3ijlRi1Y+c7msibSmWDc8bWCbYLB
FtGJtqLeQimJcNIFr/j9I0rnaNwQVTIK7pqgR0TehaWOu2JQIiOUQsWEOZ5XN7C7jFStOelgVn+b
VAgaaGviCTG+32YwM8TEpM1JvAPaAGArxdF+OV1Au02Xg9ytdOqCYiEU2yrQQpiYnIW1LY1nl93s
kHaZiONUPq1UAVUwPu9ViAVffhNsgbLuwypXL2f9TH2XkWsPQ30Yjy+aQfRLpm7UEMjnWKv/g61y
ESASnervWpmalCukYso/MCSm+EFO7TKqvuiGW9cMSkQYYpyKoQtSsQVAt9OIWeogllXvOZBI7zm4
24ssf6D/9DgLRvRtSCQgHWhzfPb0QM3caRNtcr/XJS8IiA54TkIYFHisjUqWQr4+399f7EBKaEEW
Z4R1mwtG5Wtr7/bVwDLlHNJs62O4bcCRRcXx8SqkpJnv905n8RTRCP2rQCPk0pNhiUtn+mUfNI0l
uAYbY8YCtZwnqnFsTIhgF0JaAzn+npey1iUzi8e35q/STfWE7p4wGMDnNbkb/HEVSZRvy+lmZDrH
6g71L6TjJGFzLsVxU0snCDqtb7+IDkd6hrP4dR8hWTWCJIPOnpKPlADN4hev529kPRmsKigZw4ij
GDlsG+c9nOQ/A6BtKmItV2XjNWvWhLst+DofcOpA/4SngYlx3OHYiSw1k9QAJ0GpOO6R0miWs4IB
ux9ln0f2Gzg+at2VdqEix7D8sfFGWaPqNN9Di4CqizaP+q/qphbumO/Iaabt//XizlNVz5CUCFC4
XJiAhFV9YGC9exxLSEUJrOqsrAGXPLbCvDA59mAY0yL6K8I9Q0xvHjoLhpk6H4xSjsotJvUZsiMs
cGLWHXZ7EQHzjL6U10TYrbpeXufWPP1+MslrIsnnFAWwAzKBZ+8hjdjoI8sOK8nzZUtzanfDHsl1
3IWqKy0c9fvcMvtD41c64X2voqqQGxdChUfHG5Si0RLAvOh5Va24te3it6DcsZ9lz5lotihNIZf8
QLbilUbSRpGB3ogfLWaTzy5dTdeZEmw7jn7pV7myAISLmU3yS1eXN71XDaRa/+OAHOzK9DhJKNbR
Qok3XspI00xRcgDoZ7JAGrygKIlf1nW2/3BIxBH1GVAJrcOYGJfBkNb2+tniOam+80zF4InGf63n
BkVuPWiFl59I1ucnfWJBQwpU6Ae7FDQq1eDOh8egp8hgMbQh1/9N+X0XdRSOGDpZNDZ6p3DnNQxx
s7w2XR05LucWFKwzsr42vjaV5zBkKad0L+cxv1lqb66Y2eAZ4Y67miJ/H5GmXPVL1VsfvVv6TnM7
Pg9rx67Io9V/T7pB/572+Qx6fPrZNbk79LxNG3iJhsY0k/BjDQIQkbHzfVbZydKmu/p/T2hv0wvo
rx+ZC0BkHsO2XkbIDkKqGwMf882UtiL3a2CIMNjPGofpYSRCJOnB5j4oOYjo7LV9IZ5bUajrTpdF
VUb3Q114YOfxcwDWFSgkrSKj55r/uNUNgJOCOyHe7XIzjjZdzdoU73XQ8mf3PKJ+EWYcfdAenz7N
3Brqhg9/Z+bCFmLMxP3RuM2ORHNIghOP2SGJfh5VJzfn4E+bdGH/HKLzqT56+6jaeVmm0CHmi6d/
zaKRIX5R0BnRc7XS1+R7PmJEAxiD76vi2BAjsmi/O06kgd2C/pbH7XawCI8Ao7jIL33yeIIPz+v5
AmES8cbBFDHVwfQ+vEHn4p/h3dvJPLSfxcSDeCOJx5Zw/Hh5xxf5EmF4eWZ7YWgyp1MMXpqJrE9d
vu2jV9EpH1dLwNYbdNkXMmT4ZbLsivAtR1VmDDq/okpi0fKiimyjSeW2J/XrlHjjyuryYRMwi5I1
epesg4O5aiS4Sdxv/uDDICaHrcP262izhfjW48AVcwO8rKTqdbJYejwvoph3+yY9HNWl5F7ORtMV
hy1n3aXisMSUAug4iAgqkBEsijDnGEs7Zyu48I5NtKBUQlJObI0fjAAPyP6QLebpKUv1t9XuNVe2
LWefQLqxPI/2xmGLH0hpOspusS/nMom9rRr1DLX1oX1eVrBtzZudWmkv3CEQ/6kXllVjMyCX4kuL
IfX1yb3dwCjXGhMBSsdiN9Jnw5TX5mTDd66p2L5OOxOu8y+YMsi3iThbztt4y5uYaimD8PpCJ8p8
+1fWod1vIEX0DEQ9QpV9mRYKA8Qt6O2h+G6/vtxUwA9fak+r7sv+QiWyspa02v0obALXsjANPi/l
juyMhpfZ3Txl0N8LTnJNHEd+FWY5lguXtzeDCXrmdc8m8nKMiuWkBxMXSlNBQWKwYbMhTmovhlvu
JPSiP+LeaPqGX6H0NmXHJmZJpzUe3TmawqZHM/U33/7s9kMb7hLqDDySB6fZMY5TjYMEj2FmgE79
PqI0LPSPrTVei86wGAouc7J4fuTzv22V+kLqulUHQ6w/pTH4fvfY9NVA4aV5DqzJaFyz+hKj/nq+
rDwqvtefveeEhnwkWmgpkhBlufUvW6KWPEuZEU6VJ9ZNMBi0wCevLfWTYsoTYt6lq4SP0qhh7nIt
/ZebrCqgVi+JhpnXf/SlRo3rrqsvboFQ06J1OZiemQVlOHrc47D0KgLnCtbjFr8kIaaCrcYt1RgP
/HYjkSC/g67VRxahoP+6XUMSdSu32FFzlieiOKcUp+6+p7ta/qkubkpnT/ZiPKTB0ir6szdt0KCu
F+ekI87uygEjIfeZJBW6KMpRl7ToFVbsp2/psunPnYkRpFOna9YzAJBHBt14i5OgYeLiH1xPHLri
Z7ZyueHdePlL+zrm+o7WwhLsIJFWZ9iseGZGpOaCPT+3coU1Pl5hUIHOvJA7Y7ATDm6drPHdc0xK
07/5XTaOvXPBVBgvQVtrhpbw3ri2znKvTtI5qMfn/MTvJLGOOxl1cIqZ3tSA4UMWGPIPOGUMSZ7q
SYNcLPvipC/aiAFhc6dKC8CKoYj5ldXi0htP8+49GynKRp0tY+ZIBlluAzT5gEjJPu12t+AQ+37B
GcbirGENFDiinUPEihp3XtdkhUVmPUOYnGXbEMeRB3nl1twgiv9g7YJmDCnlrtP1mUkrCIz2FZa5
aIQzUvx5j+SWG/Yh4Udeozkxf5vpC3g6RoYAE0XY5h17CNzicUb6ZbL/YcAmVtXu1mwUF4HK4ymJ
AWzOLyZuX67U7657AFZ4m/iYbp5Z1YjUApLKCM3PI3v2WgrX6eqDDho4KojtA10nBJ/pIFPrvODb
ai3Xy95JXp/55SdklQJLeQPqpQVRnjbPFUnuWGXEmFVqZCO5j8CdXz4ByBGdqRmEcL+f/PXjQSj7
Xmu68cI2jxn2UW64eUCN+ax3O0n981V6QeOrACcxfgo+ZqArzfOBCz5RmP77C3EWp10WHxp0s1gy
PodAZKE74ueuvmqWGnGUD+1L2lFAzQG9FlsffxGQghBpDSNa3L70Exwu6rkFsb5ZMCu6LWK5CFYv
XCianXfR1J7wAsvO34MVH6NEDIP2dd0+u4R9ZzJ+ECm1EuGwoKUHCZ8+QnuRxP41Rh+nt40MbKGJ
r6e3jX2/s8NsuudEBg/gN1vO1kA1sW9WaCY1hdIx3MGaEk9zPkAKxBlceJUrniOP0JTESa5NBNjH
ZiZn//ydaSJuomWmJm3/Cq99hUlm5ibczEvPa+Jvjy9Y9JTx/Ov6IY8Jmon12WU74Fu/kKK5fqJ7
tZXjM53U/oT6fLhVL4cWl+NMPtmOW1x65oDIXFICSfgUkPPFVzJkvxMBCzdzmDjp+l1IEdXEZ2Rl
AvVSQh0RaaCXYb0A5PhticMgMDLFERr0eKyvihpNXuYh245EYb2oQMlQVZZrCii7hNr8WU1ENHLP
CyKTRLTJh1TWmbvHz+pn+Wm8LSvPFzc1+pRz4IDFeEiRyGZ/TvwcPr4gjgJ+AGOwPJ3MwnZXVvlx
RVP8HXFLmiaP8xcXAVM9j2xP1GRNTO7ddBYayGeV4HZRdG0hkBe3UkNgNiZ8DBObmMCewRcT5kIo
rS5N/v6X2+tc32ZXQtE6gPUpeEgBTfXXmYXCU61CSfLmEv4dmy56947lA2lTEQXBifuOGvxDQkkp
b1cCUAxWUJlXxvXrd8dUEJn2+o7aGN/Lgrs4LkNB7+eEgufTuCcJ/Fuk8o+zNfAPmn6WtQHGiJzZ
fYNedIvnMoAxp7EDqCoh6KgpAcfK3RkqcGZOFNPHpFp9YiAA+Go9ucNIs7jOIKyw4iZbOrbsA6Jk
R6B48RAcHZfSGjJhYfyN3Y6/sWF/JNJXOcfPQ5qD/jas+fT4T0trVRrVdzjlJqdJYMt2vNb37nzf
Fk6LCelMWYvoji1f6BQ9AqWbg90tUNKJ1xluZmpNF2tizGgEz/ToT0R1ETWM6mYUO7MgiFb8Qfdy
Spf9vQfkUy2v0Tv8ev1beB2QL9Z8n6pkYdd+nNVRhFYTuQn2YQloJVHXxgVvNC1wRkOayE4dEAvK
F3XNks2OOWBm1nPvztI1gzGd8QOHACzbdCp6WYWUb9Q535wT7Ifcl+s/NsPTiRM4qF0TBHC0ERq9
VoFMoofLrPBYK4zCgTyNswcOLTEflfqK4Ui012EMX/3CdZ+GYKBW/MQ8Tv4fcgaAxHUUymJyASzC
dLHpGHb2yvl8yWs6KAlrI00tvVqTewom4vKNtgbBoWDUTNdhNIqwcpe4naGoFgQwyBf8BetJ3O5H
2BJBYlvYf1rEDBcMPaSFN7ho+gloN6mIxoE7q0yGbaLClAI3YHxokIDVRZMXGzh+cQrKEBZ5WoX8
R4ibryiCBvCNHRHIa7TjpG2Va5XJAvhiNv45qfhM4lYQLMJUP/UOv2FUBZFlhQVVaaHNuy9YhZNr
O6MWG4rFL52NuLraHeFde8rd6qxtf7fQusWDb9/8Uocm37QwkoUVfSVycXTcWK4ugCfjNdQO7NsM
UeoRp/rVnQVPSIVaGR9rO5J7Wl2jQlteVNpd8iDcd9/kXVEcwI2k4Z9knuS+znCvmI61j+8A9cv4
1K31EBFCCETpqhz2bZ24ZVDr2jMcWXMpgFo+MqiiogH/zD6r89CcKFS8yBSINmsgW3egGZ/WmecS
aeSJFeHmaB9B7y64bse0k1N+qzqz5/gUxW7ZMYAKtiLcvXrXvC54oVojCoF1aAHttMZgkLqLbp5a
Iu3VbNeQd4fI5d0XLBCvF/TGiqC3rmQomHPGz+YWHHwLt+hvgHkviW7ltuYQ+pBcUjO9d49R7yxv
pJokW7gBnxGSo/L0/dfH9SWlpFKvnoTJPU2zbHiXfOjTae6nZvIFE4HXumf67m1SsD3s0NJGJTDm
n1HL7VEdP5a0GmFB+LczBZhGZEP5ZvzMd3f2vpBbJdAsbQtMF4bwYpmjgKWE+nmIZd6m1k62Ce+e
erI6uzYK/PMmJqJUmh5yBqKk7PYRwKE0RZSYeq+gfNpjktN37F/40ql6577zOAhcjKLvHxW67W7V
4WG60gWbnt5cOW1aSBXeesa85yBcOfnqkBqZ7qHAQ93oqwdj1MsVFAUV6aqXsrrxHcWBdP/knXXK
nCyEH7lTnuCIw+/4hJWeEkmC/RDd848cVEj0aEpX1QMQUX4v9geHt0VtKAJXee5oOFBCkkX24a4t
cHuWTMCRhsPspdHb+NaSSkaV7BVNAKNiDi4F+ewGY9yjjltrKjHFDPL5vtVGDIJI8lz+B9cqznTo
RyY8g79iC4lci+xvli3vtxorRkg48fATq9e9SfkJB/psfzr9D2NAMqp+TA6qNuAHwjI5Z19QinXV
cKoTMimoY22JXgzK7klVtwDILPGgb4pWUdrQ2isWf/KYN2FRqnWeRz+8aQLPe1q/4QjnbSQD/QmP
UbUJhqRXTzAIfzPcWzZoZpgZP4JVbitrEgumwPuo0WG/dg8dPGLOZcfn9WwnBBp38a5Z5GfE5+Tq
TDAOdSlHLyevIiugaO7I2G4XI6pEP63CL4xL/++GMRP5YeAs7gnkycfUUfCHnzq3Gi2Q7ta69gNH
2vbfyWOsyQz5M3277Fwnqy1PeCLk87C608hQ27u5qX4OzAPpupw5i5CX/ZrlSbr3bY5+Sw4aY0B7
8HL1+Oi7XBUTb3a9F5nTll8z4OzKyUwC9+jOxTSEwABsRcuFlGI5VKKcGnhvFvmMPWCcwWj+NqGN
pAaDrxAHr/5k2ou9N1jDcbjtNUiNpuBuTU434zThcbDGpC/MkyQaV87n61X6bUYqNtSv/Fzv9Gmi
+8Xe9XptQ3iIa8Z22Iqka3nC33aTZ0v7UvNTeis0tv2+BpbM3+HGzYIIIHmpoovdWEu8k0YioXjr
KSUR2D7bR3GLJ2nLsKcS++u5A3eTc8c/z9CmBZh4p11EELjsqxj1CLdlkbGaWbKmDC+OHJmEGF+J
iWpVnZmP2+4QigyJi3Mr2z/s79rpikMyGOFjLmJkOIFTpNhHDMTpbKhG1gEWTyW+MdD4j4U9vuoG
Mp/JJH7Fcr5sntWDfqxRHFFW9kY+fe3NHLslmKH6r4NtvUTbRHYG29GPZgMvvkIzW5OMVRvxRiHs
C7izXufgSPoOU/3yx7GBq+iambrR5LnXzMvzoOW6cWeglzJ/7+O96P7wi5etNmVjFFNIq1AX2Fri
sue0T4ubJNwo5Ldpc0H2yxBlePfQ38Gafh/D6fK52Fz4V+2k/+wdkW7Hjydu72mI1EDtT6GQxtOs
oqrgFA+sXIFJTqnYdj7KprFQtlNJzE1uZBiybjcQ5JZSwJBCDSiTkliKONii4gISG7UaR2qNxj5X
G1P+wMx2s3J8+g3XqarUGSH7qMZu4GRtsuq3Nj2uJntgra0FNZG0XmzkQiHLya1UFceK6eu8s8ZL
/tHnZboU+lLqP7QYuc3v5kPhOOOeXshlVw5Y2Y1UWYkFerN34f7BUsfg2fzai8Muj53WF8sCVnqu
zNyVnZZqVGKWYAsHCnfMa2rdPcIeiXUS2yZYxjgWasWRUtC2aRBp/9i1+y27hZOcp0SbDjfVdmK7
hzXDa3IAtcrkcCtLnNzXV5RwpTOm+Rp5t9kTOs35bRactQsCCG9tmMHYML885C5B1afjlWUgNcKS
4A4npqMpr0JkZdgAFkKY7cZYj9v1/c56J+CBA4hIbHd0z3zQeHFAsBm1EPv15uR42lWtzH5pVZ+U
Hd/Eh+rIKM7CgdHdSi/HJbzRXbK4HkPC4T1kbA5wFL6qNUFGThPCR/cSqIae3tWnK7jgtstLustL
mHOOIf62pYP0MZc0rv7rg/C5Hi5o3ArgHs9NuOcPL5PcdROYLfeELTuuhcb0l28KNV/6JvRLya9B
0z+Kr04f6evWl75jcbxFXr9+wbpaoQiimZ5COEZmaEM2eYmbF2754Bz67M1PTAgPmL8O+KFirSeU
XNFHN6InR1Myet49NqgQ8KeTNTryfuCMQLFXtXadx4wjgk7a65RIVCONrInCL+XZ4dg1uROlAz74
MjB6TX2DBE/f3SCqIjgQLIZiS5uv+hLX5COlpRDUfyiFCjGYb+t52z9NVcJWcVjukKlE3Wthof+c
QO7EsTckVCKxZSuEdR/8DxgKI8NTx2eBcYn2yHmzWhF0slW3PbY/xq03Ka6uRwQM+t5OHfrVMWav
kAcBlXyyx4QFSy5ZzhnnbHRp3FfNuj1ApbWdKBpVtDjU2y+0mHLxVXpiAtjM0oZd1zQNqIFZW58J
vK127yBIwcsJsiqOugD9UZbjq0lI3FpcYuzluemBz6USDLhLGwV1iL4kHj0cjUsPA7cPUUVUhkfW
Q+JsjowhGxc+1tGS5LOaiAOQIRDDxgZhhLyQ0IE/sE4lb1+SrY9tT0xDf4M7I4hIc6yrJm1JUk+L
uTrDC6CVPPTKm0F2QRkHlv5X6YJ8Wie6jYSQg5C3JV6HwF6FqL0qXDYRQq/flzgPkUttoQanz3Cp
s68zQl5QQTy01pj0tC1VbxSqKANhwwVYUguQZRymXN3sGPq5aR4xsB4+7e3YqrPSjAREGl0/big1
Xr27+lgcnT9bPN7RrbMcAgD/sy360nXzmqlCDoiEUhmvy7HSm62+Nb9fPzEYyVMFaDYW9K/LS9e0
dTUExFC2ExormV4qYrSozPzGmGJ42HVYi77OFyvJa99IhF3+aCBOrOzbkyUgQsuRmEPm5Bgq4STl
P25p9EQhfnKxcf2LDYBenQuB5/WyG6qYGoF87ceJvjN52nREuCKQgDan8aHaPMzvAkZvvfQZAeKz
/CDaotlbAFgHd4UVPAZb1C60/hqFFg+4g6UzzaL/FTpTVDNgFc258ZJODW28551ItIbDmo3/RURr
HH1IkVFDtbZG11/LeF+bIkNTxOa1XGuYbMCawDuBbMZkPLP7rsfx/AQ+0slNj42VKyzdaPWIHZbv
2ZYtRV2txqTqt/rmGQQDhYWNbKG+EAnBjjKqzrp8c4pfqW8lX0xXe7NVwIqx3HJEaO03ySjDcKGS
YJj3B4HzzPZWoEy9k9rdWmjokXIDfVdwQW/5ku3IUB5c+gNr7hvdZtX5hcxrEsKq8uef+jZHeuSS
OBn+KzWOuOhfboH9zOuWhtYSls9SxSDptE1ngIFlWK/mfDMneblup51ONWimhlXa68YE2FnxVtyO
wVmogeV+wG5lOtuNlEAAV3HtBU4qucMxB4BgdVP3wB5TEIW2doEUjehvhoIA4zwN6btE48UK1dBA
o8+Zv+2xluUz04acehWhQfbAWFN7BEPobeb3Lpgw3N9IFLefH8ph5PgqmnuhwEzyZznBBJV+LF9B
6Yzm1JcE0NP3uG/MA5hy/eFxdR+1oiU+t4h3gYCrcvUtBhCSNR+SZmFV/1WRlghF12KXARBjsRmG
TBOQQ1LUp6hZ2h2Wc0Nb1UZ9k1ZGUbR8S7eLYEpZrro+3E5GVGFoScVd0AbV9EIQyQZmGcqPfXnz
ak5RUJ2DwCmxD0NkDba0c0PMudO0z3MeBlc/bJWMydhaniF/ECy3IBwqGMmu+Hiz9SLquEIhVzCR
oXTvZFo/1jYWkuFUmqk/imdVyTVvkZQIW9Iu8Ag3fFC16ZEFRlQFdBaCSUVD0ItAr8QhHucXQdes
5PUqPgwZfD68i11Tn1D1d3CphifbgnbVzSxMbgDzN1vPaTKEq0mP9Y+1q/kpYeWtL3QiS8sAj1lF
kc+KXm3EENIbSSjrmWDy9c57Ln7IsHBQgo2xV97Wf1rBllhkqL+bxwcQg5xaYT7yHg6fziutst+j
W4j2NL4HueEieLdltgMR6lllolfX01fSdJUqHpKCeqcN2t61H0xppJVoRE/gmniMIkPvL9hqbipN
b7Qs6+pgMC/1KBbvMVNedsGS4AX4xraFQIX3JXgjTjYsVoI+0CA7uvc+mD4DoSEDlsMXVqjdIkV9
YA+GinyiKGWB9ZYNFnhZ10Zw3o9PSVlkxt0YjzoZ77pjiYbI8r4nMlGfz6mCIKXnPL8bNeYRIP+w
tbF4Qz7irpVjBOFYvzW0zOBc6oyUfJ59uCE8x6F4fQK0AFHj3R596VowhePtjP3+EElFc7eWLSMu
teMZNTBj68DSQcafLt3ufJTZYEyip8jwOhn/lMlMfWfTpAG5W9osclOzNtgijG5rBZ9YcpcqQrNX
vXwzAX2QB9TiLi0K9rD9HgVFUtJuwYSqafhW0cUdmL1C6NC+IwllmyZXPhb6Kjm/6btauV3yKoNK
0PRikHLBpL/Q1xkK/61wq8dTnsBLITYV3dACGi6yKInwNf5qMmVdv5qDjAAKGgEflzYsPnK3zdWs
PKQ5MGFFFw0HUeNhIfCUkqwXZiwaTWzfmuGsOcLxcI9Mk46/RyFzl5LhQQZsVZR0q2QbDi/TeLqZ
T71L713XcAeNAd3AjTTG3wKAKhy/tK4U4w0yAzGtUnVUXa9DJOB5CE9O3k3Ddq2UBQoW0dT3V5Tu
zKMLoBjzeGJNiRhE4cxlFYbxzHE+YVhvexaa95e96ulfngEfVu3KyZs2Uvf1FjFds6BuNm6meO0W
QOBVmPcq5OcnwSLlO18eF+LmIwJWndpa3BuWUUW0Xx1SOjyLhR9krtQk96DBc1+E743BLL8yGwtZ
8Kd34sIWsYTz48mSzLdQN9p1tVcWPKxeKv4FKHscCToSGsL6834oGiYCa6V9JLiqNJKPIwkihexD
lJVqEQoOAUIsZr7mRrjw++O5fUXrklv2C9ynUeXgKycKGSyYLqCmTSf6tlxgtaepLm2QcmWe6Shc
+QwryBq9HESVvRgAdh98mLs4xYM+Lt699UzONV3ELLelTLZ29+i4S6lHYfhM9MygWwwIBdpYAMbO
Q1LoiBG8huNGGbTPGtNrM/7MqExnAiBVtL6VKrxFrsYiQqjvRO0vYSqbqrukotwVCsYp50Rh3xrr
OxmXJaZ3axmOx1gxyJMhn/CQz449kjEU7tM8YRIx4pEecZO4on63gF76GkYpHF7+7BYMLtlURWxd
uqH2FLwOMqnUih55Y/ks5BHSckmDQUdYf3pkjbI5k+09zK31TFLsYn3xPKHu54fvuWZ29JqBmN+l
R+W/WINytLwrnHHxsRY2jgL0ckvtWCGe+Iu+pdAW6dkCdG3ChANODcH9gElgJC3a6cxuRCJSrtzn
BO2juyMZ9AHpllR6vLFGwY+/YSi7xXrF7rXmONxlLyt/HhmObBizspWo7ZPuDr9iDMHRtDLC8gX5
rfNdd4Wdz5mywUgijpUfzyJdtOzYDyLm5FWheqJqnQ7VncYTu0wZ4mw/sJcinZzvQyEnN5Co8wNl
lo0Ep3aUDIeJ/YQ3hRFe4S7edxeCHkwfqbhMkkhy7Hhyb1dOZ2LQDDytitjmmAnR70IW4VIOVR1t
I+Gm3cd/DpqJRPrzt99Ln/jUJaSjIIdQqGC4SqNbxCsSCEOb7TkA4HTAYwzcX7Rk5HkfElWy/cSB
/EQeWiwe5NOLeeXWorN5u21lCAPWFjm6p5AsT187ET2qxevKDIAT6UAM99hVTUWzYAlAIv6kpGi3
yIA9xgL0EJH9o3wUBwUmQVCwpw+hh58GUbLDKhx/AD8g+b5TqV+JVvmFyhTHLZ39aQeUfYeCxnJW
RpEJlVhgQtWdUY8GO9en481sxj6nx5fGOSVA89GJmP5IbDLVK671bbK1G6Qzi8vvCNtN7XZ75BG7
2NVaST7ALP30kGS/dXm0529QabE28GPSCz6xN2hGsg4QxT2GFDI1iP+2UzcqcpNWWtenzQzC+mw0
IcBoG+eon7da+Kckj9CcMXA44+5RhKk4rvj4XmlJmfbTnOmb0e7dOO136x4V0ElQcHVrb+1bwTg8
bPUQ1dDpZ5uJJOYvXf7+2sBqt+Zr1ElZAS4NegJgiUYpTetPzPVC/B71xYe6x85NKTeVRu3fXL9u
4YyyjJsMBqSxzIukp4099pNc53SZ31XsfFNhwDKjI2qZff6VJpxWQZX1PXvMjxCOfnHvF+E/5Z5n
+W41sZ1V7Y7eUzCRv9VcQ9YUA4bh6FW9hgkwG3Zu1mrcDOtZGHIdP1fPG6QjtK/E2/2Q1XNKZ6xo
3ICCCcCngatrfEMV2JyZRQAvkQvEk4tH2lLdLtFVaIBrB06oOhkn23ohLGQil876FgNeUYrfQNZE
UH0cc0+h1pDZ6MYih2xFhkNEgbNjVfu0FVn3O2aqvFLUdaRZy+1uXt0A/j6r+Up1FHXNRq5Xtqu6
psNoc2pOcdzTSUPG/I0aRQzIcpzc9JCC+yM1sO6RjaxAk+KPL4gZfvYFSA5AC9oy8hOY1KwUpjuC
GDoETN+AP/v8kHo07t8Fbs+yUNpLGWmX3SImhWSq7/cBWn8JPaDI53CnJ4Jw28r2ALSGO5vJU7m9
MMy8k4IJMspwgGn6emX9mTcJLn1KFt94RzhIotu8+uzpbcgf7zCEmtktfKwo5sBN/xbd34utvFFz
mTw4dbf/Yp4H4sV5LrMpBUL3FvQUgJxO1P/e3BCAh20BuAcQ9x5rn7OhzHgPtLgqaP2/j1JEYCEX
/+iZd6WCjcmfM51y5VZpBlEteLw5smczKKsb0HZpGP1M8xE+udkSzrtwVHQuNnXGmkg7QXTXwLDX
msxz8Ez9bUvVwgrTdr2E3HtmWcdAFtGhWE4G1ZhC2lltWR0cZRodDRT5ReCL99c8auCuYg4Czxai
pkpOexErXzWEdQaH7yydJpfdlJmUbhShVgWkoquPETwyqUKWDgA2hbJEgF/2Pz8ItQBbeDITATbs
1rGDeXKPwNHPVt7bv/tZxpB5xY7eQJWmQ31ChW50epKzZi87GfKDSE9iXZUweDGX2cvtN90h5eS8
FP24aJLxWOBIDdKOvkiLPrxjfh/TAw8DeN3DQV/HxPX+fQueTtFN8nTC5Sicq/PBshHUndbdce1V
VmQWIogn/eY+V6oe6Z+YM5oHmwgeFLvDivvQKQOEvtxppQYGR+FU2vsTwETejDOJMSOlP7DQs1de
J9MNcThohNGXHxF8aAoPALvwTw93l5Lb0KAe/+Q8b3drj34YKE3+JdohJ22YyO05CLDTEhXiv3h/
rzVQ+LOeQ2DkQgP3QJp74+icxMGxC2fcwVUlkK+J0HZ08Q939fTPIbl8htezGr7E1vQjVd+t00ei
hCQjjxb7tYkGSGWBhv1cOJ03N7XIRCipEQ9m7agobYrx3z26a5c8suRyuCcv/gYJ1TuhNqGc/EBy
gAwGmGPv9JYFUg+iQjaFrtdRK4/AbNPmYOVjpmZIoLSWDxbcYc5VIL11aNb9EcoSaMcGJC9ld7Z9
y4Cv/gToagHjETdoXcwwtPyZ2EIHfYh3ca5nUCeSFIrr0K7cg4De0ZK1CdS8X3IiMS+tktRCZVZH
Ku1g2joH/it+VeZ3DgOLxPURMdHHXxLoO33ntdXwnqLDp2p71jI1zwVhv3TM3eE35IXvIANj1Q8k
EVpSUAdcvh241QL8XYtZqKg56Hu/cug7100ym0SAMP4uGi7TCCCXfrGJD230PZd1hiP5724g7xxy
PNGZr8DvJecfB+5CnRFr5VUVdLbOga49oLs5jumuWEDeFg7XUlkckw75xQkETNlC5jhfd+q2Qq19
8PPiuKx91PnWQoROkpZnVXduYb2VeM4sifJ3x50R4P87/c9UGrvZsu9hz3UvRqBqKQ2jMYsRURpA
LPnw0YLsuKfcMT5jbXuqyUvS3v7Y9MzGgTwHF4jshXycC27HBYDND7Dw88yWFXeUNpQAByDH1MwZ
8ont9o2lplBQq3G4aHgd7qqwQC7tNIMpxIqohlaEMLbk2TVbapCM2yS9kjuGNBLQKLZOckhKTCfb
ClVDZf6WK279BI6jCE7jLR5Eb+QwrUofM6MGNfzxQCxrJ6ENrMl49HAZ4aU3tJiyFSPFglPcjcBX
7v2P/Th+Mkn7kPGT90roeT2GPAuOQuLHQLu7H2b1mdOuuu0bQQY+vN7l8hKzWn7cioLAeMZ+p2mL
/K/XtwegO5wEZFjsh1qdYfjElqxungJq/9FIbnmeVdqOF8mLYAP/tEa0jFP2zymqplvpCHD6Tt6p
XjkPWf9Tp5Xfe+YN6TZ43qFW+jAmf/3VHqP0DnyXBabspkG32zyqDNzZ3oVFvMNT31XQKs8H61b+
Ym9SP7wa4YrhH5DTgQVs5KU+e5mMaJaKi2CPChKtnd1CNqoMmhPLU6Kba7xOe6Hr02FaGz4PyLmJ
HxyExHqhI+ckKLi3EYkk9Of7DkXC0SuBa/Lf2RWiFYIMVrzhb/max34HTfF0+hMxSIyQxUPgvVs9
nVEUQacMAK5bvOK788iCS3UFvtKBCNhdPXYKxG+nyMtPMIU/7x3U5nqFa38dJExpH0Aj3rEdt8x9
UoPEzwsNQKCQG3xHGdwvovXtG7sbtdUfoEVH2jgM9zt2JL5ocfELhVVobhz2dj/mGwNx1Sh6s3ot
NDM6+3dJECs8bIWMtN5rd308j7jZ+l4cRKCgHQ4FmxDQgzs/+dq9lOPyBkE330z/hsQ+40eUGT/u
uXJLirVCjM8WePnWG09AfJxh967j4VEi9tRscQRhMMgj9iwYwH42jLL28cTkuFfwBJWz8vx5cO9g
t6+UaBUmabdiC5VRcB35KRNYqP8UZPQDkAHVjgE0sQLfwFnJENEdBajh3bHDPdGn9bJG0ohvMA5T
38onUp5OaKJPzy/ezre3/dPmtBPUPxEuzbx9QpjxBhQpoFPr5aTmmLCZ/dOC5tU4+yKi13+h2p6D
XUKK/b9nHsjZvImZifEyENVmMu8UMNlBrZ/cKNYfq6fmnUqy4/QGj10t97cvqlkkXeLUvBJQmxhS
gpHwPDbpaLFzZHKYngPF0y91z3VU9djpXJXS7GsRm5en+0IjjlR+3Ldd0YzI3DVUNZHX5svP34nG
5SMgXeo8JDaaHIxUnoDpLeHIg8nd4L273hk5zPfvXYmExD1Z2jsLGW4L6N3LC4C4bDe3QqEitB8O
JfCI3/MlAY8wOx4QCm0dTydMW1hvEFqqdErbEwihcV4OrWHEhPeUdJ9UKPy87vMvH2Zkpct5bhs0
cVNd8tbOZ0Vx6RgkMQWMlcaBK0I27dkgnnaH7jOZK02gGat9BsV7PtAIfPpMHRqJs59XhSHbCeQx
63Xa2c6c1//eKX0F9bFrKUz9qTOTOZ0UFdmgpVBBo9Fz2HkbyvABlzR4MK9wyL2zdN5dTOJXnnTX
/9FzPECMEx3KzysBr6w49YD+upr6oRIPTMywjqXP4FoMmvZeAOeSP7p3Cnk3TZKzIgfnDlh+vnLe
tZstG4tr4hRpRRkQtZmWMYnPYA8AMHPNC0HL6pdfpZWxEs0vq8c5Zz+iSy35MWrgCTuLaL5CGo5o
/WltY6gldsMqnsqA3zS8k5d1oaKxN8C9efA5PXVPmG2JL1QqERZxSPlgC5o5WCEp9vQUAUtFjAnT
lMQUE66PsLjg83J64JDn212ALtsmima+e0V/WoYva3U7FhLgfdke5iaKW2AS36dRGBz36WWN9CXl
lZD9jZTAgHqRVRChshx7Fzuu8c/Wq3Ftn7xl9CdrjGc0cNYeSC/JB7juMxd5CMDWl/0M3hX3+fxM
FoCFDdYvGjJhNJkfzwpXj/cEeg7KnHZ0OVuCuhq/UOmMpl0N6XMOGWytUhhLCdNn65GmEfBvJyVk
jiAmxQk3aRj7P9dD/Aj2PGJAg0P5RGMBJ0SUKflugWMfm+jyD0OrAzTnxpguk8PNEt6K1JgX/294
jNj8TeEgMvLEfIZFpAnra2dlJj4Ku3H2zkB06D7TRT9txseOAXdj6EMHVzt++2wvHjGKHuMrX/Ar
phmrBPUGC8H3BIZPhqpyDGwqQAuX8YuA0lHFnyg2HO7a7KfjImim/mmO6DUpg6fel3xKtRsls//g
K531tvE2JMw9gI7VyYUjm5NVye0rCI8udVw9+7eWjUn2o+KIy6YZRKlSr/lzUN+NfvfeVzC8FbNr
Y/ke5uYjahyHD0/UJxwKVJRVb9cdHMrYy6fmXwNLuvvnvSOMCi/n42cjTHOz0E9DuabJQTbuv0+i
fP/ePENRcsrcGYEVw26IYG6yDyxNQS1hb4IK6eyxiCiG1b90aT/dkt+CdVyAGpoUZNI1nyZDJ5B3
qKrCVTU6z0R1WirDbXNTxa2XbN2UwEJuI8FQP+iXZitHjG3OzzHBzMnqjumKMqVragGhL8Q8SiaU
t5I/ltuhiGu+qW7mC7HOsFgo/SwyVmYzemSPnj/yjP+jELKSNJd+VsbHRS0OMBNcCP7cJ+fwB17e
JuKfU+L/JMAHY+HPFarG/oCRXOET54kdU58py6g7VOU5DScVjCPPA/9hZPUASOEDoubg0j3Hv59l
8S1OkDKClXkrDv2Z7NTmWEN6Yg12bqrLQfB2VZSS82qI495a7FPuSY0wDrTlQ1gV6EpB2RoZu3VT
1MFpKkcPkqUvL2InzVExU8kdyMkO9pYWb8k4bY9w7XfyRrfej0zp0K9NJgmuAjS37dxSNDEUMG9r
E9iUskEIwUmjFe9FAe5htjbtf+Z6Sig1O4pdU2O60CnkRWq/c+g3yr9FS6yWsyATyBa2L6FFF/Zv
2tIB2RY7avh7zeqdPe4jWxtbzHdhr6pC9fRt0r7v3boMsz6yu4ySJMoauCTs1KQGredJQ3d6SWgj
B9Q1ce07tlQLHfyeS4RfqInC+uRT2NtlG3w918T19YTjUI+VSIQOGZDWiXBYhL9ORkwPQ/uyrat4
WDfwWKBSisoYwghyghOQCeD597vlpIRQw8lni3gGXUMBlFLJiG3a6Jgn2YYTQsWUXv98pGhVJ3Ef
nTRUf+jb2Qj/1Qrf8ceuDKEBUPQ3Wu0MDZP1cQbrKgeW3tudTQW3gElO80+TxT6uEHrRT9h7Jfp7
CeFnY1CZ/U33uiBf6bo8M9CxTAUeRP6qxb94VtEgsmqSqedoLu59ynlYYq6ZBw/EBkQ3qeePKNCA
wCek2Q1eUgDtxFdRkpUS9xb4Vldo413KIrdjuWbG2UpL22RZX8Q1j/JRaoy+PA2yoMgDZg+SIxZk
EWs8+rmWDIJk+lifU2oz7Tu69ObzmGB/JV6s/so5MUN0ZtBLoZGsCOeiEy0hkitA9rpCnTLxqpB6
QURr0cTC3e1uzGxg/OBdQ0y92cNLlK5uDoVXpcCG/O0nYl/ei8iL6CY1KAb7qDLKM6AswXYEjxoG
7YSvsFzo0uKAyz3ylm2UeNeOxR87jKCLEkrNrq/KMpXu6zR6W0rs3jgbK0rrfCc7SBQJYw8ykdnu
g06e0afC2mdISTm7Q81+ZKe/cp9+cLzCxYe8qkrc1Xjy0beHrmZnu8QLbF5swdbndCprqkMuAhbz
JTDxpLF9pqYBNmqFQ1PJNYd1FhfGbUcJxSDV8NTi5Q2p6UFGi7wRxk19oPzi5oZsnjQdgCrA4UnJ
qzHDGQJRGKJFX+ZSEjbmGhAl+lnZtO6uHo+HwOBaxAE2waOAxUJ+KQVVOE5iV4NAJnGfnaqunELc
Tfxd/3LdZNuGLpjyn/JLZuGAKhxKv4jwLsKT/8qF+bgFusyOFtiH1MbHJ8B2QQcjpBKPU2KHs3vk
tN5CGMw+6r9bPFau7tfQjW3VAte6CkOrdixIiTd+SFrwSocnPEGWs67TwkkAji0sAuBIgEvcayrg
zvfVvuoilixQ79qqXsU5he/P1rDSG3zDz2BTngiUPs11GC4q4QbipWuBWWoWMhhPoEpyrTzAsSX9
Pkn3oqy/W2QTiFksyaQEDpsZSOXOdClLSW3n1siHQbWPdlFRii4C9XWlfMcQe/RRV7uNmmftf+Er
NzXUn48SUswuiBnn2Dy3moyMLnm1LhnFvaOZvWWvIKXKToMlEmpBeFNu/1KzFoohsRpJNNfiTok1
5ausn3R73oTextE4kWhrrPTeYUkd10TGl/ht3OQPKdaO1YnVGCdcp0QDeIHRjm/yH0XdsQ4PnuS9
mGd5wV9v5kZZw/joDZs702/Lu+qCZiOEVFxSikREh0ZIZDzBrMO+iJHZz+xgq88TY9ZARAVq7a6M
3mnOucmWvtQ2N+tZ44xcDXvcT/4a6SfOx9ktyFGw32YtDRxzDgLMQaf+zRsu0EMruFsgQgffsV0U
bdo+ri9cHMeVVeigLYDS3An7kG4844Y3Uo4HY1IeM4rysremJNvSQuhz78bP2IbD5QRdnq/QI6Bf
+RpcU/NQJEWF22YD0mi8wPe5XiD7tfS4ZnimvvxDiaTIMYU0MWGwiZ3Y6SBADmb/+8kqDcfxjqKj
DY0BTPq78Z5i/wbUKiSOn486hOkCisneNC+1Kr29nyxNCsMhOaHkzeF88wzJYzKzzU5jLrwdSaLI
6uKoyVLccpmwXB56w8cTMn30LgmvdZ+IZnEZBhR+HiJYs7LK5DrNQNIjxVQ6ytVmTeoIGN7Zc4B+
IWx7lUx/Gz8jvKQruT9bDiG9jCPYC7h8abIUH17FWhRXKC3Hmo59hlaUCAfMpPn3O4KnXWo8L3+B
K/9H1085pKRvkP12j2eNdp+ih6xlpOcSuqNqaUHxr5caiUrow5/oKwGsCxdpI01/Hebbs/O0aKYp
fURDNDakh2yuRjS/cQaTVZ30UzJAtSD75CdmslXMzXtAxda2xqpPJ92dm92nM+XX9i+FEB18/OW8
RRWQidE596AO4ufMv62I/P6B6WNpiTJJvzJdLCUfanV2vklASmZaFW2GZUlCFGJv+39UaWUw66wN
Nsd5AHgL5KRh3Fjw5UShRDw9GQxgaYjYPt9MlRpMgCulJWpAhAOw+iUM4lUfCD2FpJrmYLgQgT3R
5ucfMLOShc0UdyFKBGZiuqisFzxdMzWbRXatD9U7I1v3Tr1B1MuOuD8VeNZzIJYRuN9cmGu387x4
UN77kseqP33cJUJZrkYEDysLbLJ6gh/DGjVMDQuvmewQPRnyFAL3tg7L3m95UogR7ZYWWQzZvK7G
PTWqa2dR1oepmp2WH9JIs2HkUXE0j70Y8dFhhSXfPDCYZiz3D1CJP69oCZxogrUP0IwkXeiyDng1
MRObwu8SojXb2fvCx27HMVtW7IB3fGn/UTwJloNgKgq2QDFjV+KOx3tXtEFkk648xyYM+A7ZE8+s
gLgRMc1eQ3WqUOmWIdk6esXbxN8Ei8jCcb58Ig9oAxmPX1LF7YOFHhxuGdzayM+z/xg97/tptqJk
APpnko+FI1oY8kfTVqAPbdRrJmEMuDyFQPgY3JeYVoXjw9HdrTyOPmtBwjG0RmdVz6gQl2VjWDuU
klcVLcAVRx3tB77kScuntm0721xImacNxYi2Vsxx0P6SD7PKuSysRJtO3oP7IWIG/WvlTdUMlYVF
1V4z1SVWpGk9jtcWY9+N5bMhkr2xVWqZ1ZqqWWxjRQd/pCzeA0KvAD5RsmzKlIXXYz6wvz4cRCiy
G7C8rWg5gZdPi9JWux1p03qi9EFmR3LVn/LB8Mtd2FM3IUwe3Sq08AXG6zbdMlniWZfnbgn26mWR
YIXNUmDxf1S4xo6bMJ0RmU3tjf7xMr3R4TXs7ZI8JTRwba5Z+xaT/L/c3LjuonoJNynchzkNHjHr
0ajiV57v0eGy252CGWkISbKdG8v8phAf4/MYNlRPHfjvW4doWmTRF3HTEl9YLVp0NfbzxAAreiFA
DXXOk2xVWyK9bLaEp/Ey6rR8eJb8ZP4z8eXFwLNMdSAyJlFWSRJf8LgXshXXmGjKE10xwEX9ZZ4F
h5uO/dwFypA1vBtlASJf3WmhQohlhu/3p9HIr1CXTI2VxBr0zTP2QoqFGp+6H97vyTZ69gB5w5Ie
Q5xrznH2NtPRXZnzdO97722vBdcFgX2Yhs5VHSSeel15gmhDK/So8jX5XPpcMKEDO2RiqlqJ5M/h
cqAKdH8c80u65AFZB0HuYGWq9PbcBaP5YmpC7IsY2ekDuiHHzr+n9E7UZKJxTODWWtfmdlAWvVFM
A28AuGg9Qsn70PPWriQsltpbqBtu4OvnXxX9za5U2SF+Hi9Y0kx52/GsPKO69SdGy4fKFQjbdwy5
gRRgP6HyrmJk3Sjj+7ctrykEIRGDuljTAkLsfrMCaVUz+bdD3D9KAyaU3AwhMnRyChw372WkwNp4
KqNVrc2Lh33QzJtHragwoA681NgzXj85/1zkv0xdmseUigSPE6+NriRtNv3sPvqxIY3UaBDCMZZy
l42cN5EwGfM2UULgFxt9y5Fdj5ZYo197zdh1cSiZKtgq2trLYfkyrp6is1gaqttXQTNALmbqF1yg
wxJFYwA7Keacg15PvvkWaWLibBZDUESy6Bbz4F9j/IHLNRH/9pCLXXoU+FzuFAu2jFsSibWuCBpN
EaQ9Opsl4zCyBz6SWHr9pF0mb469rJOkiW9xj96kIA/cFnIKUkxeb4FCB+CdcC2ol6DDWONqhqPQ
BvH0mn3E+cWm/RLWpoqzioXODlE2b4/rQDhNZt34vobG3tuPSjgWh73pl7MQR0Sqeuu5bcIXftif
kKi2q7+vNNtx5SM8uY5J9n5vMNbgxb7kiUFAQVnbLeRbHx70ZsfSPMveBsrCyMvNXecdhd32Uzjd
UabS2XnUiBHpTJvp56kj4d+LRvHz5l6+M0qJQzN8QW1PJE2V3yoUohTkMFXgMhi0VsW6jp6WjZDj
BYIGb3uhTbDZGfJo7Jf2pwsDk2F88anazH7RtU13NT/QZz5mY58CBWIL/II0KvQYEwgVC92ShNtj
WKIe09QDOjnYpeIeubHaeaYuuwFmh0OpowQyAldnO2dc5zqqXduAnKKIZU3rgTPOUMGvO2IuBVFV
mf+3chkieLC4ICDe7AMLe+gAkkrg79AhBsUQrW+4vfBG99T68WbYz2aP9+GikihmMfxv06/JmUYH
4+G+AQuFD1c4Oe2Gp29ej577O+TILOFOsB7s+lGn8j+72wzLxyni+FlbRSD4seKhUZ0LH38bmmWM
jTm3hASwui6cCLamsqpxpCXmLr7Sm8BAnx6W1WzOLnFT63FR5xJRGflozwCg4MtK6MIol5RZKc9O
3F2H8/+CBe8vTkL/jntLJegv53Iy9AEQ2QNJYYq18dUDfsxGn6qYwwmvPpv5o8s1Zh5l/tiNmako
VTg4GNz0ILQoDrQG2Ngbd8g77Q+IxirIUsTXKonRCMUA/eCFrlgJH0JijzH1gHVirphdN23sa3qD
JSqGMhJWU3LY6Ht2hcG2t3CQ7icodyv/yScM7VXzeo/aRTDTPf7s5r3wouWno1u1S5uW5cuGxf2z
v9YbZAdf1RfruwolMV4Lv8GHUkWKuuY6SSMoJMK5AVhiKGSIxfK7pbiek4uy1Y99kSwXbUcWH+MY
VeIBFAE8rgCQy8o+RXcMNd6bo5CTHF/1mokkNFi0J5l3kV7bGuxJlXXe2Wtl3GRzkq6aeRIs9HPe
VMFJrsgrSg2+UjH6K075a+CNKYVDP4rt1Y1zMpYsI9hB5+mxYNsDb2Bjv/FQ+mnZWnYRTpX95thF
QVDuEFKRN6mH68ycaICHwjzP7pKnI9JFLJNkITEdzVR85IqKHy/vx4WAiSIguDBTxgYdIpFucfcE
8mnTN7Xc4b2Re8G8TN+DiwkN3KTEpmMzWMCvigGARdCt5EI7o1WPuUYIOproLiD3krJ2flviW9hG
qav1L6nNr6J81Atc+EtjhvJ8bCpgLJvQptpO8htr2OxIWk0xh8/3BG8OzyR25bhxkSaBAUP/x9OU
FROMAA5UDX58v/k5+kvyApdyY02nZcbgF9sjDkg4sb5188EshoIHBuD1CQJTf0USqVnOu3WYyCh3
t0mVWtSErsqdcfgFqbJX+CPGluAw9hgThEWj7HQyW3oWokPYi6dH0E8fPC/BaQy3cOnMNU0OmwLq
ngz3y1NtsnR+NhqZIOW2kO/tFzibIO9Bcuuc/FplovBTNlnIBCqnXh8qSl15ravvbK+e9Lx3BuVf
pYtU+qIGqP7ro1UPdWKECVjUTCLd6/7zA+MbyNorXwE56Bxh/1YSotbvQVX5/ZIOYjQufxkWAfeQ
TVELiKZ8CwI7t/rjW0UFZUXXwsbTvA0mfT9MDlfLbdzNExPtTSWcm/0RsJ0lgHYfV2DdXWBZOBhj
5Gzx/z1mR3txDjGkeqNJxPgL3Qb9VN3gqjVZCXss+K2WrQIe6brF7TVlRfvYrY9mgDQxPjqLXiJa
HeD2P/U87q6jVWExtjmqK6ltH/6WKEoWlPdNIpZeMu9ZWsHPC273fJ0RN0R6VgMhPNtelerTGHBT
4rqx7Ri/gg43F2QvuuHH53WkE7eYtrnrW+BL/bJhuZLoroaCWpTz4xR/uImgCRPsS7wO3GQ8sowr
5wSNN532hBHCJWaIwOZ4M4hUg1vr/MNKI1SlSgIxOlE+D+ZgS2oGWqY8qRc9uA0y3MyM5qxSsimV
Q7aN8zK6qnoa7gMlagD7V6rdr1wMdUS/j0+445zGGuJmYgrxREQDcLhMnv196tSML53kcNpQLTgH
5VzqNRxgQV0fUN+23VIymVMKcSBUz3pVACkgrsuFZhD3sadwr2Od8U33mdOGqwIOj+OKCh/21hGq
kDN6PEjrODwjZVpx5nfnCeBFm0XtBIDpK3k+J5o8WQLdL+DUHALA2r6k1wxfxio3VS9mALEv8iV0
KniuqU6FkSWg8ozDQZF97bn2GZJzk3y0rexM8dl1R5O1L9S439+gmPK+I82KhPp8UuSxdie9K63f
Wm/Rqhpo/2YXk3y8MPP9f4ZrhqXSQE9BpSMWT3y7U8C8iOHYVTaRA0fQbb6Cij+yP1yo6yZWB5r/
KDgSm/02c6+juFEH8i/aEIeeJMtNxzeBNvtK015gYDyjLU296XZGbsiAdRHhsmTySs4nLcP6/Qdh
+X1nFMdrMWikZ1OhHz52+3zyCGK2OR0Yvpyh2PRHESMpCiKEI2qwijvE0m33G81TlwumplcXH3QK
BeUm8OxRqrA4fQDevhXXhFCh96DoDJ7lznFtaLGPosLKZIVFx9UekHMRHvKn1Z9H95xaX91CEpjC
KVzMFCqvzc+hnclhDtRrmX1ElglKRBMORF5u21iZ/CPg247N3grE8uL6cZAQRWLHdFVPnBfzLypj
DM3TL5T8sigeeR9VBF0bafGvREg9qzTacjhYuTb80IHFY6Wka+wx2ah8K43IbzCsDbe1ntxxhOBN
bMb5+gXlugTqhUR4aQETqaNoH+3BvKVJiA2ze1Uw0M1UO/nH+hyG1aKa4RMt1evPsaRqrJo2eqDm
6guBLFRl84y6MQnglX7C5kdsQQMf2cQWED2HvC45k+bIJhuDreVs7pAQW074w7Mpu5hnmRcVn0FI
SLcfx7PyfQ0s0lhVkylWg1f7QQYY4JRoNCE3bP43VSnsXgrZb9IEnxMI2uwtqG/FNl/cYKgD7csc
Xhd/83Wd8GA0WZXqWKw5flnYrsydiqlRVScwHJECsfU2hPfn5YkM0po3T9tol9lHc0OHkylttWOP
jsHKP5z7pviD6UEt3syMrePQDlES9d0+WbJ4NozsWG3dPvdqlzuHF6oNxNHdsUCaGl22jKmYZobN
EPyuukHYyv7PtcFfUlKFOrdAfMRcGx5gzBY4EOfVaDBPYV5+a1mIEkv4lBgBfXjxhBCbzaUvPBHK
ZxXtkWT+1ilKt/w8VUwemgdb1ZWCLQd1s6nDQoAKil2/OVbzHdp7lTRrevr3zI+huYxqgTbxzK5H
WP9PZd2f6wXh1teb9r+w1V1RzrZZTk/q59erV6a/sCtavAVRJbH3GB61hQ1ca56WbdhvmCw9EDRk
ZBVp3Ly+vHFxZaEzgJtIw/oZc8VkaZfNi6x+95TVNtuf83Y+oqJmFqwBDOr9DlfaliKmIBdPdbEv
F82IQh7H6hS9VvDEpyG7brxxk35zXPf1ggAlJq9O8PpyLXPrINmyRe84zJnNAat+mfCMbroh+3mX
24pJGgCgoKfbFvjfoNynXchqfKVhA1OareR9tNjEe/rGj458pGYMjLZfR5yXnitlBVuf1lW3AKIh
YWKfGOcCDH0Ab5EyGIoqQAef4A7+rTQUwhvpuzH0kxi1+L4vhCLBSCC31rA/sT/B29WmrxY73qSZ
RBCQBmN5upESlmefoKq24a5kJWoJkSs61+uAd6ZYRWsTRcMBgK29ZYpYI6GP4BJPlnfSgjprY2DY
SCSiGoQUFzC/JyYyOvpOqIMZGuhRCI/n3oFCXQ/19WZLgGb1Ed1BVv6/bXV4HWkh4eEwdazQmH/T
Eu1MFFtswpxbAlJAEgGQTUIRxi9LxGxxBa9HWYnz+zYD2XPfZvGo/f11OhRekJZTB8bLiprIS6TQ
aZb9h/JR+mrxg+q7hvn5DiLngNXoF6y5dJ+dnfkML1fmmQf7Tjr2lGAboucQmpGsxIbGhqbjfSoG
1oyW5S9kEg4bPm2SHhzLIKu1byaavjGr74H0jK2eNmeK9q+6+XE66n4tLd9GxJ8VLZWXobbcBnHH
qqvI8OiefPLmRA76AIWiNOVEoRXyjyvns/8OlJnt5eSg4nE2z2ppZTcgEQ3o5k4iK4X4838W62dr
4MTSdbYEWdlh3ey/NrbHWBMjbtJNO31Xy+lYoC0hmpn04oNtEVfyXj/QgeVtpG9nmsSVs1TeJVSQ
TucYdrfHet+d8a07TWUPiNHWWfw2+IxLnQi+3kz9Tc/n63BCZ49INlKAejuca+xr28hAxWJC+Bqi
tf5yW2No/v8bdBLi9oE2XvE2yW4JrDVUY/V17OhxslAx5cBjkk1zvzbyJftYvfA1biv3SOLNm2D4
PB4M5oJ+Kzln7Rg6/L6FWPjJbpgryIEJVKfVivuTMedYpLhBnGLYPtZNtL/jGrLH6TcmZY7egBQD
qhpGb8eo5yXEukdIXmPRsCdmHqaTrH/bp1a/cm2JEym8mmNPfqDR7awpeoNvKLVyokO7BbMaIjg0
gHxTFO3uStOYKwbGAvKCCl+pVcstOpjEhuWtQqjbdJdHhO8GNo6dFsz7yuA3u8NNTKu2O0rpZCxk
wYqZnFIKgYsZUAjr5JmzyhZs9PYl9SHqLkDJvJE8HOBQHZlEs+theSPTZ0K2WPhMcWpfdfApC4QQ
OL9qNGs/+jUMb2r4CNxBNW9BTw26E75wVJzgbEvcV96hf9INTpce5GRfiIS4htpHhhG65pDUZJJF
PQKCs+wTxKM7VddhivupcLfgmK6tZr1qkpEVf0gBpujkwoLWn8xr5NLxswNfkxAfiaIdV42p45MN
/ZozQCLNw1gsj0xF0I1+LZHss0XG1OUmchsBu/SUhZMrImmfQI94WrAc1ZVOaKyutC7z+bEI79gr
d81d/Hyl2t67aFBrLDCySDfeYpjiqxBfrDEqkvP8FL7VcJOK+oHqiywhrCy6KgJXw/GopQKEvsZx
aJursS4/jHtVUf427bXyZyfOG/uoa7tfRNE7MLu9EusY41wV++Nh8yRYFsqeXXho8sDTdZiv9GVT
xQ8wVvKCGAC7fd+lRt+50KJGLLdkgNWQk3hyjuhklTdwNfE2yTwCPzX2OLCrKzTQI+cWp+pDDIkK
E6Tw8OKSZ6w2iIDfuOegQADqLEMlTy+x/+/KrUcGhCHb1T74qN9SfCQpNGlk+jBI/Mbcmq1sjqx/
DpmK4qjToE/geegfRZGRj4TE0vfZlt0xKJZHpTcPJI1bTWbaTGnto8kDbCVg0M5UzidEkfKnV482
01W40PwIqeaHet2PrFl2jbxIE19sXZmObOHj53vE74va5Xo14iVBk/QYotDrKfefgqXGb/BtZRD6
mM4mkk1BJyZFav+h9l0bscN2K6bpFU4TRi/dYT5TR3KBWoHX4Xa2zYnr9njD8hU2InTLGqub1Qi3
Zv/HPdvfBB07UiBoyG0vxNrlr9bibzrSGHud/I9ciJMOrBVLupxDnlCaB6szBBSyxEQK+rOyvfS9
ziSTCJrlgjPPHsY7n5kuzMZ2V8+Cw07WXl08SabO+kQBgDjwvvAWOBvLPL9vi7oyxhNOLh+H4FAs
M9X3dAidVMKneYKI4yuRjLg4s3CtH97wyuzjXUDs5+xXIZSZfonKvYx+f0WeqGfxdculq6YL3Dhe
JbExSrR0efZp/LfcTWuEwveupEqRzleN1U5l1LasIshYiS/XkHCpkHOCy9HOzSRHEfrDO4cycd4E
rq24BGujA0iZ0sk39opjMq40yfycD6bXEML4GiUD76wOnHNoxkYrWgpDJSSZ8Aw67sTF5fmfqg6W
QGfFl0Te/YQxVVSKIhPD/KqRFAqD4bqZU7YBzK7wAPNCAikTYX4LQNIUSMtBQELTO4FJM2OU7Xkx
eFYF4jfJGW98IOZPaFX3I97reIXKLgrercuvoVnqWQpS/Qp9gAmbdCwb9A95BGInz8zrzomRs4VT
Zh9r0NKZldrwaZmzcijPDyz6MBmH1UnUkaztjrZInsmKS7NiBwVQ48m/JjLzpKLRY19CAUJGeX72
EyenOJVfAIEMpaPdxC2s/3PmDJ20uf0+mQxQNSFKyX3Q0/+BzdZX87Ma0CXhUadnNFYSqPhbukWJ
DNlYAQqsek9kWm7Y05jtMsKIH3Q4oKqUxm0+xuDNSbetox3EtIx4xVdtoqeckJ0wT1ccwqgDs/Dn
HGKh0TI1JV5Kltho5cy51A0Hnp7kLTAsvS4732LjaCeP07mwJODJb5ySBC+pQMOrNT0zRXNTrVJ0
L4Ziqy5aggPePeZPttpQLrIpkWCwJbsKZsdTrMi3xEiyxi6JM34k4Mhg3qSGEDtfxOMlFLP5AAXJ
UOAK/RG1t2iMfHqW0TkFrolJuKyKcZYX13dS6wZfD7ZVG/dh0jsX32lt4OijTR0kBLO5f3XrT5h6
0VjUW+q5zlfW/3hIhOnzqzHzFLMKGDnsjgS31AUdEJovKu8g6alcfxi3ym41ekXurMUor7e9Rlhw
IMRfh5Owai6Vv2zNaxgJly8d60sDMn4pzaNX4jaB4TvKVTX/GiuKjt7AwGi7h2CmBLY51aokQINA
fcBPhs2njx/Qm5tRFgcs0xIurYJpsmEhGJOUyWdYbwHShDQfE5GYr9+7ysZae8275qPUt9Pcp6b9
njLcCt97pwBF1MiKL0UD/SCglQyaa+6KraVDcv8kRPPSu9jacGrYlad6l2sQf+Pb8YmHuOBUB2W9
L3HO8I8GohezXculVFuimGh3UF1zeN0nsn+7UpZhGdukYVk/LVp45ZscP5IDtYSY+1Z0HlOupcPa
F6YsMzoEHDELBYAK02X+Q/d18hZcM0J4wlVOq8SQXCizQJBM8XDLfChhAKtFzIZMOURmsOdVsC/q
XWK0QnQZ2emhG2R5Ug0bV6KFt6AufJ8m0vBj3nI1D0T6SSTAOpNXVzyaMmjgVMmKKd9U3pK0SizV
P09PnkuoROvPjZTpev4oAY7prsE2ALi6vbmdyC7eSgla/dxNHG7tKv0Mr6ZRMNYzHNCWcp2T4C+d
t/V2a0sEuut8N+5VO0SeL6FtwAPCpXnMjGyurz7HqwlAvSlfIF/ImOpyedx+NgPZ4Hz6VWxIQ01B
dIRcPvxoDyOXCS0BFahBCfRR9JyGez9ipkOZ5Z8k0KI62DzNA0+8Qg171SCv6imsHZUhlE0TFgF1
b3ybsR5HGySEiRBVw/kM8uHbEV6ewuxj8q/g0ULRZbDmaTxD/ZbjrtrAMeYKWDv7OOy4EQe+OLhZ
wjBpXuB1gWYZXTwi12YqHIX0kKC8Y0AfMpT4LWFE04Jc3tlExTovk6IPcE0sgF5AqQubnwAJ1l3J
XtorpHt4WViwDVMcHkVwuUI6oTIDmfySiVj2rY/way6wyVHVtI5qPxqIXbUpcYwIq7fU3sM69uDe
/8XY3VzHwPHBh6IUKt+840k4Fk5Pg69X02EWiGW7Zhg3VYi6EvZfQn96rt19aC7qmTn/RRQi+rhm
7MzQ4ovqX4O0sE1Ysril7E/nBb5KvRzez2irc9DKfKr0zZnlQqGABS73ZtCBt+RQcS/TVkFjMhVQ
PUNcHxHag/c0n8feYyQClFbEpDsPvPwOto5zJRVdqZ8FrGM7Zv4sFd7+ibLoFFTNW6nqJKJd8zgH
O0nqkW4N6IMrKpvDXpqsqNtqNUl0I6Aq2RumSEFaiLfQaN1h05jVOBM/w8pABVUxuwZafwWDVkef
dXkLWfTOtT/FkDBbDySjbsKpC3UZzPCuF/opuU+N6oK12zhD3lEOu08Ev24gKomP6aijaeJW2iAc
/MCKDd0RuvmfhNo6/1EjIJPO0sw2aaDFmVqvUfvXbOn/UepeX75zW1NrQ7sj5S0o1dvjgY3zncll
ZjX1hSGfkp6DEqDDkx4ijDB6YMch/WqaB3uMGSPm0fDjuySHG4LWDxWndFJXNE6HwDwTtwrQ/qyl
1UdqR6Zi5Xe4gF7LhxqZBXPz4QPUygDaqniOM0bVxxsR1DnEemaXAixXLoSAbtfiY29rkeHaH/Sj
jWOazWG223gVRcTQwpbsA7T5rslDoTQdLNVx4z80eu7Kmokc+pUQaLyrStWSyk5mBJFUoMQ15sHR
Mx2fWTprwXIQeb7PhUQrjOxEDFaywg58p3HaVSEw11jF/sEayH2TfGDLAe5ALINauozZi606tTdt
vd464QkfVwkV8oQTTmqelT3lC7wsOqeQ5eMKQKFv2vU2Q7a6ukIffQ49go7Esy06HfpcV/YTjfoq
N6j28ezXX6HMxDp4OiZ2v5mjqsADa/YlU74etRAC5uhKQy0N4/egoK3pegifRsuc/f95wODds9z6
a8ixrYf7MSsGWsVID61hehmoo+ht/Kpv9Ts1i5P5A1SFUvY4qzlL0uzRW8ziG68+4EsG6xFGTkYw
X9PUMhEZ9fNNoYz/JjEmrN1CB19WNuNCShQ8X2FKW2LoF0xbDMLn0alGqGSwBzwlTj/QnNczPPeO
p9qHX5cxrJgq4LrMkJcJF32iATb7ctetid9MtrcIabt84cO+poPTTeb+KIP1HQLmPXQ9J5lWdJIH
yMjV7pD8IdqqLsWieGAIXK71QSaTvk2OPJqp0qYOGxpblL60OQdpgEb3hwGGFGuzLaGymuewnWfW
3pDJaN7FQ4OomAT/cJVtpulvga4DOg+JclKUhUAGCXQ/gkDr/6nWQT5yX4ppEcmxhvXXXbXYbMyu
iQ77qJ8zZZQs+sXb+4k8TlsRY7/RWeYphoqW8Wwu1unB1atMNO3DKNEoDxSMS+8uuAabIS0h30zL
GaT1ffCVRSc3O97T2uxFWCQvVDrpgVBpdnmyB8RzvfaTxHpfrwt7ucLPW+joPE/3z+n9vRrFne92
h4znTMpLRJMSU18ngR8R1Z52cgV7HeJkhia6hmRTK+jWUHTd0orptt4e80vdiFGmabPHxzZgjRNf
h+BV8cG6HACQDzLNvwOCeqYvLS9RD8yXw3iNwsy06TXTnsvzMUmeZ84WbJoxbZr47D7Dj0VqwopM
HxI7PFNbOHwkiVexyDSKIvINAtLMw37o1dp/5IO1GHikLnuOBcos1AKUg9tlIL3oh5sIq6XktjjA
7ephqHJZhvkR13LOh8/PTItq22LPEHyuAerEgxjs4re+up7+po/B4QvngFhM0XrlH/migKbVEThv
TZqTm+rCIHjWSTBGVzjLZ/2PZqzhP6U4+eA68ZOk40xg1R29KG6X6uvSe7VoGAZ/y2kUgVh8NN16
kMNcVDxfA11ULdnX+a/yOfjZrtwUt6fOq9ipoR/paZo+TIYm4MPt9GY8Maey20cE4IC96Pfpcga8
GBkz5uXfj6G22TYzFKPU1+S3olfGxqsw1wJHTKrUFVumgtmioQdxqOKD+TjYzVnQ+K+1pDrjc4m2
HpEIoPItTjo1GGIvl5mJ+Cgu9hsFQUujSbeH2DXfM8Cg2tOOl12aLZjI/uJ7Zi/vUq9uwm8IiFQM
71t6+lAJLYsYI3s1UZHdXp3W0/rm7qxx0SL2N4bgX45SHnWmPUQNIFvqk+pfgL0dDTf2pPPt1833
chFtJvKpL7khITv7S1V1c17QW/dSlEr8PSrjSccfNrZCc+Xylu7oo1k653F/KufpMUp42ir040+S
4BAVFddeNb196bRWJJhPURO9yd3upgsTn/0zIczUjlGAJHDRRWt2t/8GWt7K2xy8vo314tToDAGa
lPCMHqYsfGqBJWZJM0RK7mdfoxENBpq4ZfeWPFv1ocbVNZ8xfYYbGKxe+evRfG5Ret1F4+ZZY8aj
Tr+DJqU+RbyWrkjcuMov4+CZqAm2e7YOd6n1zoTsj/c7O8Oj/P3zgtyt4E79Qho+5Fpx/LKz3a2j
sO65k7nvIyD7j97LCNvB0yqZKjlkuMoX0mgwhCKw7Dl9P8vCNxcd2PPlvlXsZovqBuPqTxDvAoCg
CklfGE/kVhUAxmyX9B+FGeh0voiFUGRDwNDBG/LJNRjC9m2Css2Kjisx8vBihQ70AkTQ+cSrYV5S
0O7nig8p8jxFMw7GY0lXnfd86vCfyrxIc73WvWkSze/5zf+50vASSpD6EHDAODMqPGhkTRfkJfwx
HKa74Bva6W4ckuV+sPUmj0k0xi2LQ9gfabnFgTli/SXUmpoaGdhgUrq37qf6znN2o4s/2sFfc2Su
Iv5mt+kqeR+Br9dbALkMiZIi3RNhoC0RdDO46N9ETqaKPqi4VPzgllQQ+htxLQS1IJBdazURJuSO
3oDxGxi527xSF8TBEnYmgB0qUK0J6YbMkuQ7IAJztiWj8OJ/HI96vceeAa80VkScM0Y8+wZexi0P
1rf7xm32eE7N6EwaH1XooZv3H7ab4rVDJR3zhtaCu1SOZ0Lpq7YsvGTBt4c8EVVHqlKEmloYk+N+
OiAGG6V0siedNvKrn7K9fWLj5ErA1Vqw+3bnJwIxLtGQxb9FwzrQd0S5MSrQrl3I+OnFeIa9i1TL
YQTN0oM1F5yviQQO27SJdTL2W4LuOWP+ZkRf8nQwTapoWMxo0Zc3u10XJDPKYSyyy7fIpTEUaZeU
BoVPOP0UZKf5rCAqdSIgwrhZ/cD3ozHy1NsMbEO8/PUoD25nLOMJHVj3k5rog9tT0NFLr3o16uEa
qfOmrKVJCcV7g09yI8vaW8UP5ZotgiFNjxWPwExWXAh6quGfL7r+WjSoSKpM1KM1gZ927R+wt1Qc
UholNS8mtFpIVxCuOtnf9u9oWNXfJe0Hydp+kYenEuG/ykMWZogcCkeXPXQ5Onl5iwhFZFhW+8KJ
Tezqwkj6Nfai+m51riH/cVJ9/K2SECjwekokchb4bqMtmRf0ZYsfBOMz93nV1SrlFWrNmLJU/VRl
k3BR5MqF4KY/ydmVJGh4A8UO5jl+crFUOr0RZjTdze0AaUIZ9zKU/b4ZA6wKGAAPyiqHLhDYDpPR
e8WuXMBC8MVJ7FDsXs4NtNiJk3SkatCP4CpHcocB30BCtyGqXkf/VvABSIxKL4QOuFOBTI+aDkeJ
9Aiwh5tIGb0kjWbOeIG4ffziO5pmQc8+i5tylfAJKn2HGMZNyyqA2Kv7xfNqw4DlXyIpJEeQ0q5S
7sGlZ5G6wQH6ZXvE16/tjwlxvK+WDaKaLozyxU7nfusds/UlbQccoKeSIzfi8d6B+n7UBSY5k0Kl
PlUnUzor+Jp1qmrx8wyCGZQLzrNEPQBf7PF2Yr+njPJUrwa5eNlNw7Pc86Xu5LDWwc5z8MOF87JU
r2x6WuKdsSVjmBjkioLwMvPnknB6nsLMaEhKy+dCa4qjeHyEqEUSHRWLTOlStC9JfMP8L5Y646+x
ms7tEvKTe5gwYcYr092b5hDCsqjV3w5CdvXp1596Shz5uFT/SmdjFmqf86TZXRMtYT9RbAWaPjQ6
ksFKmio+QondXoldjAVGo47e7mC8fQFyyXMdbex5figGK5lU0XQKYgs6iYwEbfT+2ddlkeH92E6Y
74L3UIN+KjJW4R7LqVUbHz5Bed9UuWjmZSjli/lBmZuYcAbM1VJQY6Ka470Ay6XkJz9KNjIn6q9n
L64bfig0hp59yU2H0aD4t9AIm6gv10Up7SP9QEEHmQjVaMNsAhr7VLgwuTVf18qS9chEW9KIyu2a
BONfC9mBLAlNn4O6deUAIdQmOMbHWFXRlo/tI8TiuUk+DdA9Fe+XAmIP6M7oSUB/DW+PzzXqBgeo
9DXiy7dWSRUFHOdCDMG6wGvuA1MdZHf45mC7fvrnmRtfmHWBsWmLfMUJtwFA3i6DWU4gbyBVN/Ai
97cJ0SVDjY0Yt2sKFgmglmdJz/G18YZwSbEFjjUWIS8ajnH5ACFCWqJFGV0D9ADoT+aKAy0MLNPC
T+dFZTPwuOWiwnJlggkq71dxFGV5bxn0UFK0uRqM1QPHC46gv6gNvdi1tWg4oZhPWYWBMGFlcVjY
GAFu+fXc2ivT2zuoU1TkK8HRKChiOD3g6U7iugrL7St/Tw0gOAXflOZAHIuUHuzkNC3nuf7cBWVV
9r96qY3umlS14x697AU+o1G8Cj7YXf0ZCDoTqK/ELFdQPtKMKQdSLqW2CFWoMqufbIMByLl7Rx1m
2NUaKEtq7UNpwKyRn3qn6JQ+J2XY3kYWkhZRk321lHqZVmlfSyO4HqgjiiPax3vplSIIcLs3bhkq
PV5umcylQ4+ZAA+oA0axeiuwtulJGnWLVmRnzUGTFsGzbVTz+yOxPKupf3jpz0fDMBKCpqHmSvtC
iDyceyW+t0sALxufg3hcRd6M2hApIwgQyycv6S50atDy8fmsIJ5hHemu5jAHip0bup3ypyhCO79r
Q7j1Ehpqbw9Hpuqw6EzQPEoyzWHiXw2A1c6oglt/1D0d6TNg5NARdHe7cOD2l/nQ68yRLGDR63bD
8mn+9Sy2U2r0lh8DOyuNjH83bQc4pgkqXXH39JYM5WaOkZ4lhfNLuDkCGqTybNaewE1OG2xH7Nge
z4zBjdaUgBa/RT6kSeEdM2BBF1sLxgjH/3VZLKpkGvUp2nSBWmV2RPJNOZosjhgFzOvb+bDx4/Sk
kJy6lrVLTg6OHRVNP9JCUpsdehWI5Iqc1FwDey0CQ+Ega/kB6NOKKi7v2m8T9NMWcjdMFrRU8BQc
FlK4B6/MDeGMjXflbpLiu9r+3CYet9buRVFkCRWSfXZoVtXe0DlezwjlOWjgQYhUtdUDd6rX08YU
9tfQLmcd+oxc6GpuamW9Hwu2MUML0xDLohbBxF5FxVun+WN6+LfgC6DxbF9xB2jV+WAipeILahlJ
WiHRcdNzT12SNpWa55Q6fzWrobktdwnKUj8eZR3h+CeoyLglgXzYs6/jKuSGyPLZQKbJaav3O37O
++QtOCQtFU7uEPRICmcdsVhZEu3vLrY6MXb+kE1CrY972cMfk8uvmRUVDuxBd4RD9irNsiHv6b4Z
T/XMANs+fEU3TirXbeKtHpV3PW4HRMT05Q4NWX1X0nnkWqFRHH2i28fCBZZcQvHaX9XEI0cZXV1i
aX6YEodEAuq/ZFFoZAvIRUrxEp5o6q+KYQT4uWf+m0Sm2RZ0FAmC4PWdHOrT1TCZHisv3h3edz6p
gUgzU8Eg6ijULibM/Mmj4DaS5DWqhO9NMuJINYQngtn3c2VIxEZh2z1XML3vdboAX1JYSAS4gsWA
M8Iv7zQi1Lzw6/dujylGLLjgqmmYdhV8vzbYlQvMgkxWZAQ2JRn7SjKDowfu47YMLhYRXH/d1+ey
dz/MrSXYbViZVP2Goox71l6kCgo2ixvRwJ8lMnHjb8rGf73g7uf0eQsiZzo19SRbLSCEEcrhB4oA
o5nYJHBuPgifAil/v6g2Ag2YptTgOlKPcpkRE9fnXXFgPtbWZSg9QC4sAByNUsLMa11tXCeyJPbR
crMjUxM+vk2fry62lleRQCHt/3DCcJOCysTaZxa32MGfOHx1IczvSFsmd4ZCh04ILou2MNaNc8zA
wANVUIqKBLSP9J9fHkJF6Nhq2MW1hh047CKiVR7Zh1Mpu+ClTXMIzFgHmFHozQgvFdEuZKmVFd8L
NE7Jjvy0e306MTBvBaBDZoWpMMYo6rBgv6kT6uOC/VcONzUCsNHLKvOPlO+OwAJyWbbH+Dxfbn6p
o0u6mpCXxv1+EKefpdpJ+Alu71Is1cPIIaQgBojqPJN/jNdrNi/7aDtv2NILDNgxjS8q4ozCnDZy
LRWESGcjdp+aPqVLXFTaf1NwYotd5cnmTETXA1fEsHn6UdM9c99L07apW8jHb3Eis/GhpbF5iYtq
tzKS7uYcpaoWdItfBCF9jMnLD9EOZU40P3ff4yGwdo1FjakCM4HF5s3NSK06q7+gPHelXHETYOiy
TbnH5csGSpQL8ug2D1kK30aJOyi48uH6ojWOYXb12Z1+ve6LjvmLw8oeiLRDL62R+0MVvmfICsSI
RlKKsg2oajeSJQNj+NuK29ZIDTKc1m7K3lzkIFFXo0qPCcEGYbeoAhS8GTqyWxNQhf0KRRCY8WOT
fNZeB80yxnwaQwFC6+e2JRjWphZYHm36TvW/uRn6Ho9JelQMJxlzTn6aGvkJtUtx4zxJyKOgl6nu
Sjbc+1DXkh6+Kv5eCHWp2nu6Q+0aof49MDIscEkie1AvDW0LbE3hX32NJ9Bac4D8ra2YrQrthx4k
ehbuQLK8RtMDAklpHeQbcm7RUNv4dXnhHpVHgE50ibJGKvo4swJECVLN1e6E4Z//uNoWoMjO/kKn
x/wy7NZgEWaqk+yiyBD3OoxtcsmNv5Rvfub1lsDy465nzmbhKmW2Z/KKdQQEjvZDEKBf0aZ3hxav
/550bF2tf1oKQKnUrLZ1ddnsb+ewHZy7MCZQRFge4OO8vHIe6D2Gz2as44jtGz4FHPUrqI6tD0de
Bn/BMrH/KjkAjPnzLea5b8dXR2JP5vptTvdT1OIw0w4XdYiD1j4joVXXmW3nvWY/JPlMDvzv3aPV
o9m9GqI31UNjIuyLFDABsehewW99NZmLrX5x+IF6oLmKQjCFN+Vj9y28/LaSEoNykxmPYHmUFxSn
nQNPu9QBmog0ehiUyNwR2+5wfeP+OpSnijtnU1BynoHz/J+A27syDWhG+oUZJlRGyhyHw0ux22LS
GidpPAEmfgK5TbeXJTs0g7eYlU//db7ZhLFqnxfIfTYlkW3qIs5yxznfAaZ2Bu3AC5IJMi+HUkU6
geda4auQUcuzHmQvdCxjY1kEyiekbYlTBsur1G1te5H+7Qgsr7UF5xtTdHBNuvgHvgOEY7MnQkSw
rXbvp7athsWa6gBVl0OQzKgMiAeKRAW2oyTIzrUc7CqL60M0DQEzvGPmsV5l0YezFlvBhKve7mgf
c/SmTET4g4PAJRnW3yWcQjiXrrbAnN00rKtM+4UMP0/lWr5+D9tVtFp98qliWEpC0NziJWH3jqLo
XDZMFra1DdtUbAYF8W9xfEzSU0e1FVzevo7hyifqU3JDTXMEWd2z/iDJ5c7oZqjjYK+SdP95Nhis
bvY3Kw0unXqn+LcXgF5NVo5ooMUtmF29IBYctk8+BRZz0Gi0aLVeZVEjlt+iCZsNjVKCRVq6MXe5
gqI4SO9n4jWPqZVjcbK7dFcfqiCG9dcrC9BlWhS00r99fqI4BfjcPp+tT5HlHsIMcslvGWwkVPHJ
E+6tWajiJCK3v8kOR3Xeaz3hQ/v4kxTB5jDHmaxwGQqCgC1pA1Dnh+Bc+MImmXBKAXu+UQlX+m6s
VVyaFsLeYWj0iZQVPAykE56IYdJd8KoVSoMr9smxKaJuJRo6XWlw3fZgIhVxXf8ns8qrOV8zSej1
9ypsudfRmSSgc/6ldmR3h4tuWYJbL13jebyKHILOJGam/jYnwxnZbdIT1TkvEZpPBU1T2oLjixE3
u6jkR+L9ItKQUXyMCi0zSstXEcalpfs06lLR6iXo2RIQjl23cNqM/szjQYTx0c462MVLkn4J9+Ea
XU5MgvORUCiGqwecDOddMe6+8lmzbj3artveyrTWbINmahUp+jg3mdPGD9ZuELvJPWfEkdV2ys1a
fCjwCrCprGUdT7aIutDV3YoaCnn/nUv1i60/9yzoSha9pPosfKlKnnle8FY+ESnCFkW+hx+27oyF
JngV1g8tpysbpjWhS7ZMTtaKx7yON8ZnJba53BGLPoIU2H/9U5W+xBB2/gRi646styjQhQ5ZL931
WLY0Cj3ZHRWX5fiZAWApL2uwP2OGEdwR6Ci1NgGQvMKF3RFR1d/adZtoHtiphhOu6I0+9UlaEs1N
hvPcLEtjf4f3mOy1Q+OPcV/udi84TgQpdr71pWBtKoxyXBzCpI/9uO4teUkgQUME2ZUkwVl0EfeJ
WUqIVzISv8adr7Xs3ZBHwxlO5mNA+sCyR8RII3hfcp8f2KE6lvg7re/IImBD7Dmhd3b4p/X9sQGj
X/FFOvc1VRBng+BVLRUw0FjwvihzVHpEeNDo9XdBjDivSJk4yEt4hTlJa7Y9QO1uxVLuB7YK/BUb
Y+2I8XULCZ10rIeAs9iVKlFW1gZ+kpewHNfqpPyOP1Vp3Am8NyR2/x5ejr7e3fwOl++UkgjxzHCJ
KNyJhgaFuummCy0lvGUTgvNSodlGqlK/dg7AJab9AnbH+HV0NIuyq1VL7QXaR+hOwJ5ZjG5XMK7X
Gb/vJlqRlCgg/LQY3NYel6Dmvq8VjAzlwrO4BukOYRtB37a32HHNxyaE13LqQci5UDRr6pfAbFHt
K2WI0hX+EkNwPTw2eURVE/gmsYaBZTVSxDpGW5yTAIIglDDnq6lUZSMXzPi3yUVwSGOfK0SPXSiF
bKmDcvvUdQsfz0RVMGf0CS7xMKabYEhvSW6ExBPh8sl+/+VqTNbOT3Cal7VVgdZdpkI1AauUMGDT
a2B9omIIEXWEnIW3yilIjixsDKJedFrvLKnQAKqqaz4KVrAVyex5xifRjMVcSVOdklJMGT+rPvp3
6dv5p0WwixxGxAt3e5yp2wyLfi1rRQY0Jo/UCJBGDALfcBxlSNY7XuPHA490aQI9zIRaB6iduF49
a/rimHHWpYgJ3KiPCBj8qm8gmSzb7NO3u1KIX9P3Rs/31LJ/5XS++mI9WMn+mfu4IRSUfdW/i3zs
sPUTfg3P/PocCws+JQH8QnIsGfCe5lU1LfgvuzSi2PdNDCttZebtyX6WgzpNZ8QeoJcKIH2Suu1Y
X+gbLZFx5D8PvRlidPZE+BzyqdIVVLHNnugCIlzLaSZvBKuVTa+BbhZp/xKP83TmiplkQBXjFKRo
+4U7hEDzCROur2YH1Ou4YvFG+d3AF0wHfAJTBMqyMYyHwClxVOexOs98EGHHouJCMblXDVUY2OeY
1jMqok1KG5hqb6A3fc3sd4XKLLLJVfKQi9Sry7VcQu40vIE6S00MOz6cfRdUPBtKNLpYI9J91D0u
7qelX1lwTif2HU0aMbjL4otBqKpf5TQQiuvQH5Hdt73BORLBOjU/ul8KdxAKr6YNaJZjKKWwHjEH
t+/Je3jvmd37q1vUtd8j+/+5WBpIro08gWev+ZJJca1FlG0oxGsFAoCsJoLIoA/c8FjxMQqUEonH
Ed+lDRkOovc1YooqG8xG9Us1sITb0QfOfHuanIWumtEMht/PaR5WYZoFSEom7TMF+H+TMe8OKf02
iTvpxjQaessvTaNOAHL63tNlou+NjJFznf1uCZjvtNmqDyse17NACNvcl9EB62tp5Pi2tmYCiCi6
PO3QqX+2HKZ3iKwAS/UPFM6J/ZggT6o2dOldS2ThKrqPJosy33Vk+CWVWE3T5J97TEt773KMosOe
MK7mOvdeOrgT9e4bLBmhkpiNw+VvyUtbpeJzlYwQefadgEXeqFPtX8421pvu7i2LGM8SZI0r7n/o
y7hz1Kw6BABjyMPIOhz0uwJNwWC/7ryyN2wXOBhslXVXMAIqCwBoa1xT3nJw1Pi6GZ/VFRsi1OYR
5sKubIpDCR1MTj/1t43z0UbhUnGgcWq2dEi/YBM4xm6uPTyTEEwAt7LTjVzM98S+bK/KM8mYTd0N
CaBj+19aRPIjVp2t7uV8y7YLXZxsTV7NpF0tui736noGDOrJMScmPdgmwbFO3DV/KUkGcfxx//RD
G1Q+roMdWLh3DY+v22htVBGzD5ohmHT6h8RDeeh66Fg4qwC0SLfmrSdZZ8f4OdKJefi1YHWsOJwU
8xBlQRupiggK9DOQ/OBzTMRmXmdg1u4PHFlKDGSR2E/QnqrknJpTK/TTyCIcnruWIwZ5z3AiRI3u
CRHogkvNnB4QgHA50GZ+HtrHrMILlN1J4o16WeQbUtUG56suQ9JTUYGjjhen2tCKvNkUghwfY6K6
WetpqQhSCqTCBhyDYP/a9/smfNYdCh5Xad6KPY9LghZ/Op7pzpOYhYDQIYuGlhs58NKdrDhdG+PI
A6x8Zh3U123WdyTcSNaoAw+Ok47LOBFQdCbvd9THG1XES3C8qzlfwc2XbxPtr3He4FHcjUDKgG6b
HBRouGWEU10E6k6h0g5s9z0Gi+ppRp0qrMv4vhPgsvA+DC6Aw4gQJcIrZvLJUrX+sTw0rPY8Mn++
o5g2HtUbvDr5xYiOBxY+4GN0L2Wnvy1QjlR7OSOKyPnfpXIEaijXJEKClof+zv4LYLg2gyOl9z1w
lD7+3rkzzkbUdXKwrJujHxWwww1ZGKXwcxQEnC1V9OonOhffoiuMuwwD3NVdl+aKXsvFZf7ogJUq
LkSKA10p823wqbrp2NXipVHIxjz2piHB2tLiBIKslednOhO6X2HL1n1l6A/M01zyVfxB3KWm+ns/
mcx8v+OyKyF7p+LgFktNuFJ5KPyYwEGzaRLlZTpKCIJDcQXfJGHUtvSf6Zw5W0Dx5n4lkhieMgZz
Ip8fKwhP9uSNbrdPnKpv9T0bMeahMgA592J80xXZNCjPH9lnlDRDpVWcal7awOFrR9qJCcaZHSyw
21Ugjm7oglITEouZyaG8siwfUviFTL93JzjljuXErCzzFxDHkdzAfO52IUTJiFGSL506ssddv+NH
4q2KtsV5fb8sD/s/Xi5PI9MJCvF/VWoaP2PXp/yHVg7weIMO9vPOG31b5sNGFllAXaQO5OgCtN3t
z6t6fuB/9gzMGs83N9Qegen+CyTDxB6mRWO7lZNM7Ufxkyk1R+FpBgNgY/T3Ql59wbWYquzKkrNK
Q/JF9vVuCJugIAHED53CakJ6exmvHB8DiIbu6/crvyx1Sy0YcxMN4XgOql+VPIyq6KFtgvzvo1Qj
K2tIeL/Jf98j4HZNwScfROZXD8C0LDxrSrKZ8n2pt1KQNQwoiryDemgIssSry69rhWSYQUUo6MfR
ilI+kjRt1b8mE1DLixyMi2/v5QOrqJtFxqKuR3Xo5yJjnI54O0HRDkQCBtXb/lJ+3XQLTDxF4n3U
iHM6MR3/Zrp6WrC5KbnOZiswvKq1hP32VP8/LMn5Qyv199pIAszkJmXjtqXBPr0fXGdBKlnhgbIQ
afaUDTszVMzwSspveXykUrixZHXr5pBatyAxYpaFrBQuJ9xaCQ/z7MQRJdk116oYmkfYH1uoiJGJ
ixIVCG9AtwJE++lKo7qkjomkyHoMk9D87feEUoXGfc4iZIV8yaWOfI6fuA+uEqvZAtPKw7ehmm2a
0Y4iQEv6M+YJWmi41of5o4aj896h3I5R2xcqdAOnOvL1rcr7zuEt45F1H33xiRpxIvqa1/ogwJV6
S4BlJ3xx+dvW0xhMRGiEGOwKqsuxWN8jlJwQwtxequLcgju1AjJSRN5TKCU+5fy5vjEYeF6UPmFW
4P/An+sufzFRYwK/FbEwA+wqRnzmd32cXrUwMOHMz/OZZXfQwGpgtKkIkb6kOq0jCPOwRrrA3Uw3
CDyFPo/39G9407qljKzj25v8JTxXiMiLV6eaoGqHXjxil69ayNI/5r65SoBCT0sUfNP3G0SN0qgj
YeN4hHLLQDNslUR0iOH+ucePnhGKGmOqKXQFtLSlHA13ZFJl9pnBAS3rj26MsvYnOZMLBYBzBD6P
AfIZqHb/BOh6+k8LQ+6BH5CJOsII4xoU1eE6RvpJ9bzbX6sGUpE46nGjbfc72190jefZk7qDxfOi
awmBCw+IqbaGpNi6I7M90hbbnr1Fm2sOx/qjR7SZV+ArAGZ76+VfAwdKTwu73x3352q9Rec6Mr1N
jXtVqk9fVj6Kdo3RF8KGmZH+EJjrzoRf9DoPTOeod3iXAzU4zjaWN25I3Y0Xu+r4Kin3yiYCpfJ7
M3E5r3R+mo3krILFTpN2rhJDC9YZehVO7fN5beHnbZUbzdMRZct5idm2d5FtdcJyIBedZXmRF25X
rzvsPgBywfLf8lv8KDtNNwtugVYhE6xM0QdnSlpG53wAjo93zVIz/uDSk+wL79pezT2gkXDJeYVb
r2SaLYUAcom5l4U40OYACcfnTIeYoj0VKHJdJYQnF+faQpAFkHIU5BeDqLpKyasr6w25BaGTKNUm
3PGbYsqQr8M3n7oIsLU4qCcZjl6KTprXP6gMFO4khZoFhocdKyV+BJUj1AuWKGtKYeFhCZvgYYwx
J1kFSTXKtmg+rWajSgiAaam3c21GmrHZeWs2A2d/JCwHslZnBA5FdoJWa5jqzQy4oVGhvDDq6/WH
hZSrxa2h5EhyY4xVFgIgcDSumAOAANxbNcq1xX8MgsfyorWd9cFOMV3mkeRk0TPCbCRhGYg9xy6D
qHVYwuqTabVjNHorLpIQsaMIphKSu0p3bQBXiVLLxhnwctVvX09/iqHc5NBIeZw8lqerdb82p7H5
Z+wP2izG4MFQQmHh2Gw1eAXP/Q/dKB2ESauVYrmAiSoZfvOjR7egWF/m3uAT/M1rgPJQfv6zpmhv
xVtYN83djWDI5pfspmwThX3RGbLYMyi3Nc2ho8Bp4q2smrN0NZ7ZjBOy1sPCdXEILVeMJimu+IHn
NTnqJ4oAOeiio5npRIshO29zmjVCeikF/nLRTN9XSzZDhoUqFhytncYpT5ebf5eA1ZGRx6CahhxL
2RcCu3V7GUZ5RYW7dxFfpvBYIeqFetb0EGHtU7aag3857VJaISeoIqPCkVYjaY4mAj834NjmRWw4
IP+FUXXKyPWhAxweyqeqYCTyjY0s5xG0xghX3Ee8ucxyBl9vMmL8c+72VGe4+qtJP+s8Bdn2Nng9
XtSFXRcs2KaMCFo3POTqSRWhxHqlMx6vW9xCo4oqpH69CkLqYYGdGvRprjbHi4ULszjdyHoCp+iw
QRzzPZYk80sSE7TlfGAyYk+EImbdg0a855kIFP1XCEr8xxOpMoFLAjYhpHHK+GJAwBVuvyGLJCI7
58IHEmygwvsitH6ypL8umPxnzIYHnqa4835ZjHh6mrlM4zPzObylnQYrK7pczZewQPGRSxiOJ5jX
8G2fXrLVXRarKyR/qKNmpR85NyqIst8huvI6GDlq1dINR002wj0pPoXAbIzFuso/auAU93CNzwcC
Wb0SXPZQE++4x5XP6l6z71FN+roXLfb88u+a1fUTG1Iq6lkpBedv0KIzM/oZ8mB6ajzaks0OdGon
PWUQAUDeVn8lPzN1eP0NTPnhtabwYJ6FzB51032hLKJvFHZK8kmoItwdlzp4doJ8P2yNBjqNTl8n
3OiE9oeDRpAIBeeo0svgagZ1KOZTRCKLVKtNHmnbj2Hdkt0TV/DjT9CF7YstJ8/p7ryW8clasOmM
/C4MQfq6P+na6cPsVVqPt1nGS8t6czIhnTXgDtYITy2rfQ7opdEgWDuxFnu4UeND2KakcOIxM98l
tX5vr7ula5s4KaUsn6mt0QUymzJBKh5J9eK7Fsqa0tSWaVWrfUFrDKhZdaZnSZ5VnBBvvrd4yzB7
ZUoqqNFQfcKN2yYsjKikQZGsUcf5R7uQ2XqvsCtIR2DiZUMrPL5/ZNoJW0Sn5yR7TrVraePWpbAi
8SL/Z4MD+cBQbnfKDh+04jdNmzwst6lmcPEuO4RJHQ4Eg546JcS4RuF8JadQ/8jRorARoR+I4ish
HHNRrIBfgXaXjYdkiRbLOrGfAgTXYkbyY6PDNuN/ZoLg5a4GAlkaWqGRWNJtmpsyJ8zi1g82fulK
+uia09wVuIH1PhjKnA8yM/cBMxUhSiYpGzo6MlJnrxUjrK0Be0a2GEvdgi9+xgySTCKXRQGhGhwt
Vi84sP9jFhcJBL4AVoB4XhktmYxc+LO/h5R5iaUlBo3MDgomIo0Je/GN9csOg70BQaqbdprcJqX6
sKqwtiU/p2cm6vdWA1bXlj27lVGls91aIiaztJtRhRBi4NhLdn1vKOdvacLx2kAKDKMNTa8vvjrM
jhr5mi1X5i75VU2r1jDWzScokqhC7bka0yIadGGEZQZmskXYUp62vwEm6be/bWEngJ9NnwgvEAiN
snGjFgZ56Zq1animiUnAGgv3mARKkm0HA32+xQM/s/zZkOUMUuiJ1K+pFjwKFvJYQ4Xjz3l4MNWH
bi1P7NHYFXlezmZMugcsAQl33BpXSxnRFcKejlKVI1WsmM/DKP7Bn5qATzMkKPKXxBbOL5dJcGVX
G9GN8+1dpcWrobdPhjd/Oe3JZUQpMmhwUT7rX6yIWND1n8HJApR7hqywFRMmLApZ3QV8Gv8QlMV3
wVgFZuxb2k2Y+jiOuhvPNsZ31wxzvaw2y2lsbAXifAu1QEBnFt6IiM+92Udk19z1tT37waDdWkxc
89RCxeH7+Qe8wAnblWYCfI0mQtdSc+oWRWTh0bmwDBtXC0ThGrFfAewZXzkUSJsxuB5rjmBWxiCz
LFiKIgCWryWZ9KdvwM2+b9MqC+gYWEMSNqbMwEWCTGtuJZezaD/npJqQMf5mU5ZRLhKw6U2W4egQ
Lk+Uxko6GHibP2JUU0hsWFOkfqX1SbXWYK0BtP9HuMzYipgqL4D9Y7FSABTgtuwPkxyA3zogjH35
jNRGqC26lzcYaDLB64YGsW8kZsyRbFLXdj6W1mH3lXZM68ZBiklpVc6QZJdfRo14b8o65M3E9Z7R
ijalQwxtV7RryU6O1C5ZrNvhNB7dv220HX2R0MB+nWpvouoOsHzXZgo2O1k642xRO6g4NCu8C+td
+C/pGxc7Z4Z04RN1EYLnMgOLgT57Nik6Itg+/1V/2CiW/Sl3hxxIs3/P4q8bqH+MXgeo9e2K8dBh
ZQwuC0oSh5Rfwi4NEmUEQdiJuv3YYkhz7m2fwtU6OQWxg+J+AYjy+/25PnUwlzg0UM4ojWwcVQ9G
OZB0um1x3sIE6sJtT2nMIJFPVeolxRA17ZGV/D/MjE+XxrUkyGIhbUemEQf7FK5dSVSkE2obBVco
uqeVRZ3s7NxrncXheqmfpg8KUKgmIPg+t7kQWPCSqP7ALdOPmFDP7ORq94QgX6SyDLNjmWpnARTg
Cg9ROlBsCe7lX5AnJ0qU7JdrVwOisolMdtL6GR5Ug/pDIlUqtKVfpopAzftEyP4WNeh9ixKsuFQ+
CH5Uhz7unVPUNx7SAlSycyzWsBVfkWvbsU4fiGg+mSIQlk9dJst+8q193lUWri+ekk+eJ/Iy3WXd
Am8S58XRFI2AZferIbFQdpvXh9Z1LUYg0nU/nxpacAQTGg8UPv1k8BxlqW3kz1vlfIWQhldBN+4H
LdjqK9LZ6q1LRDfqtrrgj397U5mJD1Fyr83WQrKif8wNOtXYHRbOEpKegEejGzGXA6AkZbRYR/Ix
Oi41RXJPxEgA7oGyUB3p0iABKL5TalwLf3sVZptJ6CBUojRohERUWRaCqiHpPlmQKxqPv7HnqcsJ
zyEetuq35VD6jbyBQPUsn9+M8ZXKrEP7MayJule/56JIb8XXs9SHqs2u76pYZtjoFhp25uCYlicY
KgjuldI68a82085tqMow02G3iTkQX2jGSbXLWZZ0AHM2En0Y3fhVctblnZSueNEGmq635hB5+rv4
S2G1BjeGyMWuJj3J2MWEWdSr1NhScSxw5m+j8msYW3TSq+EvxOhNgFdtAFGTxkH3nh/ngeBPzJPG
WQeGWH2qGoh9r77FzkNo2s8Cz/ld0GkgnpTC4MJFZw7Qg90I5lQji3hkUYvhN7K4Fe4kB4g3xqvT
r4TS70Mo9shYL7g8L5r+UFySpCdJQoiseY83+3XQOEhasz5FWJpEjOq/zKo/4Qynv3Qhb45pd8HT
BhE13dsJCAJk5t/NMnMd9857ncsrtwwzpBZXCtmiR3yYRgjSVrDWXsTal+M35IW32s/+zekPnqcy
uC00p/7DAG4qs0LM33kE8nJQ2/qiNEsJTygiKpkLclHU8BNzuFwH7+Xb16Rq3V9iLCabA5eDh/YL
RKxmTGiNxzsFx9LsvPB7s17zeDZ9Z/0+KRg9hMqsu/1PYNJi4lTxy62NaE5k4SnAP+RTIp8I9xjH
hgXGF1jYW0eE4kwQRxWu2iGFm78zWwQPC5byi+uQIMMx9whx1/QAsGVViWwLsb/ZwL3db92gkmWW
c1ezAFsYF4CxIWKGvt2jffMecoalXMZz4TtI6d3/CTrrKedIyPc5/hKhLSyyBHl0quUZHjdnAlci
mL5LJwGDTCYzsYqK/NfL4Ce73v+XmDCkSScz/X7p+o8891Di3CuVHDKBA75HSaASV6p7m7uBJksb
ogj11JAHYHCsrN4BTCyzmSbAlkAxFxzWsKcTse7Gw0R2rtc9JmU8ANqDZ4bSHrc3kOHfmvJ04yf1
NCCyyGcXJNDByOHNHwjyW2fojEhu4R4yWt+jnonSFt486gM0FTppsIGHK7m8qmisjXlH22GhMlYV
xNnCvri0k0wpplIGaLuTdWGH2OSFWlqD6Ea1cOvXE1Uos2VoRUg6p7ZejFQQK+fjiG7qv1/YeRrO
XNZg1qNQruDHjkFOOf6IfdSCh+97l4iZD7aOQXX1O3d/LJS+rxS/3BQ/EnYRQUkj8Y38e/bc18n4
8GM7buP2Syr7RQ5VBVJsjmjsrhkwUk04YBdMyAS/oP8SFRMjcnhGSZRoHVgPMyL9oHn5KktBxVp2
yaI8JLYlIRxm9zx0OidrwKeDPZZFJb8IsU/U/3445IK8sGAaFznmLGf+5RwZvssbPA7rxRiKmDIs
wzn226FIz9g9to2mpk3+i7k6GXrFc9w0953MsmiX+eFt0lR3EQvCEoevmIrRJWq822Snj4rasNtU
xYLj6HWrRKbs3mmPnENMdrt1qshvtDQDu2scAkLcZ7ZcZ8FHeS45CClouUx6CXZf4o+XTozvBkct
uY9ZWiwfug7OyxTSNWfmvwUBHB6fWiej+lSI7D/Dw27PCHTkNI+pUwPsFtVdssuC0UQzASCCFV7e
YaLCZTrRrXVVghayc7nzLP7CBWmG6G0kdFex5QeoWVF3PJtbVS2khqzjgQ7N1PYcrZB2wxaKThq3
dkrA4jHYKPScfHdUkkc8j9zxDHfF/PMTDyGkqsIzHSgfmKedGBYUDhvHVqpSd9MeJkeucmlmRddZ
C4Rrcf7SWao803O8MMrNo+N3KyVP7m+fuuZ9dWJ5Rde6/yROKihjTMPbFyRlTuAdi5YaJu/4D8dn
Bg6vQP9yrxWzA/30p19yCEgbDZJqBtnQuse9GH2OI3PtxAAq4TlI+A8g0RgB56aDhtw4XUp2SlkJ
n3QJ77ubWRGu6W+vITYMIS5ypkRLee5gtC3aVHpTeow1ozlGdS/THf5NKkl52ne6pO1Akn4jgtbe
kk9KCDPw8Kd18uzuGruFnFAFerjSzD+Z4QuI5bHEGxFQVtFuizIu/uQR6r3MldzmzA71I55596OX
Jq+HbAsNeyMWIC5tkcYHE3a9/tyqrBmbTAbSNttzR/NYFpscDHXbWQIEKDOIiyCTKXMiiwhr9CeA
0dbLpflb/tq/iiDBOmp4jbw+Z/hZr6Iw7SNfB94Sku2T98tJ2l60sUqQx0N+qAjpBtN4bS3Ln7/i
PP4jM5EmdrVBloga6xGRYEpCDRIUPkv+WOzmgYOJxD7zLQNW0o2gspZG1uIz3uUBurpU8RqbvCck
slA/5LWpZsaxEu2axRQ8gM2fEDPe6DLCOJALD/0h5mLjeMSpHNYYh7ITqGDayKv2JxiQWc5d54UR
usCZzfvEigqIGjhrDGjZYBX0mKm94YaytfhO93XcuCBi1btOGzj6Z/4YGeOokqMOp489yapkHoFr
C0EZ+z612ha7yNxKxHW8kiSIelc79gFLIzIu+gJVyIS6iuszlU+BtYH/vJCyaEH7hCwZGw0mRDiZ
MhNDRwwnl46PtKGSwWk9c5qr3PTZGl+gJwllwI57DYYNLcEGDCnd0KBF0OrFi+cX1U+EvUZ8gAlT
xoyS/dCnzR3uTLnviVpwfD7hsU06eC/Ve6a9xPzsGa3isoBjPJ7BLtP+15rNNKQeHT0E/6KLWYo9
fFdvdm+X7A7Y7fhJ1ogbPsxqcABTmSOr4UWQSLqFQhxtzBKc6ySjqX2mXhLuBSAfSNJfsxBWfD0G
fiFrX0HDa0I7e/EcwqI9Iu/YmAEzO8V3je+QUsebyrzhms9M9TuNyZrtXWOrTzaB4+EvKx0bS2+R
7QlCNkB/9CzgmPAUUUKADUf310VW8nB1K3PQi9PNrua9e8BaQfq7fgsMAczUAigmzhdMMVLkGd6u
IqAscWk06SzbArUioajnR5FO3gLF1d6KxNMMYtAoOfoKAUlcb/7K7xn8FLOgje3oaAj6Pgp+1X0F
n4H50dGyhPcc6cCUgn0aeuhzIc5FYEvjfFYqdKQCN/ZZWPEa7Idz2d2rwkaRhkffR8DIvI6AfYNZ
vcEE2v+dFeDCpm69vSQazsnAMDSPAbrVMoqQajrTSbyPg/W4r8ptvU8RxZuEcA06dI06RPhy3Yp7
td9IMg/ZrlFaCaaw5QB5mBe6H/n+7wLU63c67yJ8cUoxtAYVgwBgejBmhoMNa4n3FHKuGcE/9f8X
CVgoHm4IJQWuOj2Uz/2zQFRhgSu0TbPs2sRC4RdC9JlrlHaQchEpqtYfzPmi/BonYy0TMHN6iq0P
ZCrGgsBwgdvjgA2pVndDsovIQDqfjSpS8aelRaSAEyizzcpTw35e9Kz2/Rqgh1fTPWUSDy+ZMqGQ
SUIYycNK/CQHhQVJ5bffEA//ZTakydCqQy27yTd6M9RZjaDpy+PiuZ3u0/d40qke1CxsxjQXk04i
OHyy643/0O+Fn0ViQoGYp9lx8qwKCrVzk0E9Uwr9eIYIlJ6ZJEBVTLRaGiL7xYTqKPpGvL7oWLNG
3Lly8pKo1zpkfgpFNPDuw26op1uoO1HlzDiL6rVEtuDP4EbKtnAPwODKE3ZJkDhKusMhxFeU2/NM
nOj5h7mgtSa1t2dvn+kD6mJFGlof52wAkUjvO2jaPryY22pxB3Gjs0t8ZfZEyItRxqbYB2fmIp9p
YcTA1rOdJS9uN9VFrWODuThunEUU8JKI2Yfm4aonmG/QSsM4/iKIw0oxsVBiox+PclSkT2ebbjzM
jRo55T0MEPA9m1D+k4JensZpXKLB9tlLLkWy8FXDhBH+vBqW/igmkLMwepewQQjOe6BgNa1XlGQN
b7cAqswPWQLTNUJlAA5qDdrbcO0d4cFynlfNaZF8A5nu2YWcUhk5eooLiFpcHJufhFz8E9Xld+n8
jz8Eq8DpIJZgGrhmitaCKRc5AVTaKw2lTWpl1PXJMPPqVW54it0H5O9uCgkxzQOvxizqgc4WFgES
NWijc/XwK+e3nl00jIsgxgr24r5E9rH3+kBJNMcF+oEH/vHzmFXBjK2mUSDbsEcP6rkDj8SNeufQ
yJL4ZI4k967YUCN/lLcjTFUA84HSFYlZ249ElJzSe6itM2B2CJy6pr/xg6eBBHZ3Ng9+JD1CJtUw
Etq7DHTn73h8ezzWD40mdL9BYvOrIPr12OdKGQYY0H9d7dJNBVAYqyu0UL/JXILw6uhbr8dSxlDr
1+HMJi5PXZFrX056OluDiGqlF0pbsTXNe+vTn2+h/sSQJASb6zELMjkd5A9E+ak1Nu3/V7dGJi7W
lzlroMyP/pEQY/YrtRciLfJgHHEjH/hncNMc/mbqGDsIJf6BMOTKp8zH296fUQieroS7XTcJDEFs
IbsiNWEXYGfMOko1CNIYENRS3baXYZif833sZJhLxlnhoEtG0rH7wyPJMIGRv8vc7Pby7IMS3vYy
dvVDwp+uqsj12/iZf6hk92GfvzGUEuzxwPs6tEeM7FPnzBCsbBcFxysHmbnwKxnj65YJ6VoZmTtE
nvtqZsIIRPsDMKbc2Gd4KTGHbXQmIY5iIDPNtsohyrjINa29w2AOHRo3u4THoG7qzbk7kN08ArME
qkiVKGyCUs0zEI1eyqtWU0pVWZd/ME0POVQHqoCqXTVaA1qBftUIt1LOX82d2kMYJ35ijb9BSCGZ
AaQh7s8y1QpFkqiiNX4uwlV0lATRwbGUfrzK6CNyYPHsk9FHuxy8tH4LJrpSI2vK89RZDTSZoEEp
4B6mrO+UkeFkBqObhgu12BM9KDuB5XREwD5rYFpi6H4k2O2YDMxm2YkE+5VD/92AMMmHwZyCW17X
8wPxNYxrbM177wks2BYRYaHomg9Xb/gaz7M2DituGxfOtfIlY1XEbHb8ZRdt7r/MJpagrjkoVsDw
M+iPyIseihsqr9GRDRzYIVXMizHfb1/ezhVwesk5+v4VgkpDHGk6xBxcae2y0BDNwXQfWf4RRTLD
59D4j+3o/Zq2T+vrBlMhukzQLNdscoxQ8lQiiobeZLEMLI4hCZIHSrSi7Ue5rKPBf6IC+mTWyD9K
fJJeZ/QjxBhwPDBlzj6pOYvIXRCLw7v8+uA6rKznOsLMnTcfD4O98buNXPhPNbxAGtXayI0tiB5U
2Ropltaqy0r5A7bv0q0ZxypFGMagLwjKy9Xx4g06MDKP4OoFOuuwnohZkl7hyV+zmKcrCWe8wGy7
zRLBkwQ6A9J6IzMfCezU92KO+yElMMwu8/7C2HRe29vy9NfHhzTZZhi/RgLLE9Vyr93a94yzxawT
JIdZT44p8eBUwQpH6NtnEcHoMJmPVhfL64fyoaYBcdmiflxu+zx0SAZlh1wgQMQLhByvdq1zPsNS
50Wj+crbxItbQW53frgX50CSquOc/iCfsAcSct7xTK1hY3IpmRotEXVZm55N09GT8D030NpLAZfu
RPQS7sxcLLBw6cvEW4N8N1oGP0idXPyfW3bTGj+56czJN73B6+ZtHXOE4EZ8o52Rjyl1Wj87Hn+A
xmxQuWZpwFT+Y51klRKGjojz17UyEuYrAnvZeTYTL493wWmpprmykgCXPLLTR/8etM9HNdDTVJfy
r/2d451M0xL0kTk8rPk4CRtXNqA0R/LRAs6VMcVU4XRYT6J7A13dA/DatpwLMbm8tf7y4FmqJLoO
R89N3BIZ/OmMe+w6SLMz29RRtXBurV15Gs1PHiYitJdivPAZ/GQBaL88wN+OIi8LqIYwAtDrPIc1
ywI1136FvN0W2i+P4o6LaLuOn1VFagdwMtARRlCUtcX5jIoUDsehZ0yCokqafH8XwJ5CiGD4oyYq
AwLPAuUifflAB40tohnoWc6fux8uDANTftqhK+cm5G7mj4IgrGTn7ICKX5H7Vr4wZ1/zMHBYtY2G
8oYtHYuxPPsBqI4Mw5z2AB6fDlEWlyBi5Ioi/Ut1rssta0+xZGN0uBZvR4TAIL+vTCJoxjPAiwqx
3Y7qoDX7WJ+8YNE2B755wuKAEeukMrQqSMZoVhJHRK7VXjmLBAY5NvqkAT0k7+CBPGgc2IJlAsnX
C9RLYhlo3T42iOqzBCy2E5Gs6qWW60tUB13PEyDrBFYvSj4PpPRMxNiwlZoNBv+6o2EGZ3tRqGB3
a7cSgFTbpEPs02JsKOWz1uYQ/UfvxaAHeEcWBxSuRvFaQzOJwqp3oyVS1VSMD+4woTYFxk9g4Dyb
ZpM1F3gKlO1WvAq+BRDDEqpQOcGH9Flw45NM/Yky1+0RBwotw4E7QfQoW7q+6mbj6lhUEPLZre42
8YdGteDawuN2o0GnA8hZA0KLfnSxPgpXFfAg0qpHe1C78gnMPNqrgJDvFaf3aRITBQtW0aJ8UHan
uu+smesgwg64zE54v3v6XwdLL8iYlSKvqiDNH5JBkTie73DjbxsFhoXxAMTITSLzXpxL82fVtzr2
ZzFdAWRTsSF1O8MvbXa0FD5/Kmi3SjaoanuL67yN4ielmsorI9kHW7lGD5TpEnn87PBXwqFD1sQh
ZVvi0wa2cJ3lSuZufLdV+dlzVcuhEkzGAdyjdbFA2l5gU1zeFYMDaLssxcdOQVGvFMeqmpAVx4nF
WDY/1z3uWCcMXh6mINJwNjLnCZd9I0afruNwvnF/6CNLVJ3gYJnvG4D8v3sh0f81r3TgG3r/LPbf
KuNWGAM84Kr6hZcQnZ2nwnk964xdbn5bavY1avc6FjE1X4WKW9R3vd7eVKx6YRd3G2mV1m8kYrJm
w9bc7cps6V/L6BKqg+F57htnnVqWBOvnUfUVwCxbtpQ2UcRtlAytyFrdIkFn0UfOKfaWkpZjAQc5
apzNzC3rgfGsfzCXqCCUTFG0epqbHZhqr6QvIcRhLZCiK3NFCyGlOXdNTFYuRsj/6LzqiZxitXHm
2twOOMGpdcIB+TQ/8j8DM1BCMLhB+hka2zk5dN7iZoSWoe+2/QIuEUVBjq5iwYq4LG8FbcPIXT/J
8nJNHO3aMn6NnIOHV4QioeLRXV23k7ApIKselIydnjUvFLpbKPArUROAk+x+i0gbTFhoP0sOagIP
l4SaZgcLXFtQmqIABZ+aZDaI75dHgCnaNsNufzRFwkJtl4Y659cGdv1/yzhU8m90BPBoLW5ODyaZ
Bv7+RdSxEdEXIYsa/on+v8QKzoWqIb38z/J1MmaLM3QHBH0N01mAzdnjrTvsEsPKmyuUBhbIswZE
/ydmYBeyJDkUquBFVVBX084RM9bRJjFtL9YXoSVm5g3T1nSTeaEeUoTHWcnTav01pWFaVpOyHWRN
+cZKMe8YhwBmADXqlxu2C937FmxXnPcp+iDYgnxik5DgLiGyTe3wJCT2d7UoOPeMne1cw8JuAKww
SmkpM1EvVwHo5aMxJImhG3oXLSi7oApy9CkKyn/PSmsEIC+3vcfRPEuG9u1GTiGsVSqaUuU4ee9/
MwO1TnFsCsuif+t6W9RtY1Xsi1UGaavAfkRElTFZmQ2yx6Y7OuW4CWGPuZMX9j079onsFLlGRnpE
MoFoTrCcaHkrxoIDZOeoGUQ6hLoME6Hx8Yz+Tw+vGsYLD15IbVgVCooWhOCEsCxBcUXmHfEoBrJC
1ejwGrx3Zs8LTTXjvExdx391oiBXhRRCvujrXEYT5hRt7W3MBBBrb6x552MnAWUo4aRa5WHPW6lt
HV3OyiM2sTtufGpCKW/YWxk3fA6AaiBOamxKeelcRDmNMKQVZN9nm0/BWPPoWTaNr2LX+d1WolPD
pGVBoQg9thnFQYz1y6P+JLbNC74fkRzF70KD1MgQD1ZAXBatKUXJxzx46uutKAQhob2keOX1nY6D
TcVxqE+JSyLAsQVwdFtvDX8FFSfiZ0FrP0UMfsKBGxsuA1RK40jT9ADtWWt1nli49U0SNiLjVFy8
fFvq+Ob6yOYDG7RjENff23224VDa0CoH7ylsDKT4hTL4sOGVvwhcM/MoAXWBO1Oe1+W2p6ldgpD6
qCEkIlgmiTgeJfB7l7TjVAs+ULy3u1ufeeF/K+7Dh4wsBKNeieW+PxAvWUxWsc7JDMi3KO3imMWN
3KZxDt3/UHdPM2GIOoUEJyfbLs2oIEv1joFxjvwu3xB6hUsi4qN/8sTYV3NcxDAxrzEgyj63N3oC
mGM4fMw/BaeIju8o9opAGp9fHSxccZ7alVjDGJwi1/SZDdMyferM0uKSSm8zkewwcg4tkfkw/j1I
E2LuG8KD+F5wWuOFtTeGMPDhXN6NNZQR8Yf+orz4Mtfbv3cEd9GXsGxNpFt2QRo5ohiZLtNWEnwD
/VY25GSlseIs0sx9Xf560VqEMLdas8bt9EAKCSdDeAHouIFcFdpboCGdiZoEeUdaEQT9sJ4asEJr
BAwOBVm0bgLal3Hk+qgFvM0CeK62cOI9KA3RxQGjlwLp2GwnauJAk8obIjBLM8pDHPA+OaxGo6TS
xzh4tu0aMc7rUxHTvfbzWCKUW6A2cFHlBDmkHMa0e+h8ad99dI2hO3x//l/Cs/nuFXBI7bZ0U9E/
ZUdq3ZgZj1ytIEYtCR+wWrboRszGCac2s6Hl8I7Zxk1vmj1PwdS7jwGuwMS0E0SIrvU1dYBqilOH
XNKdhgmWPS/oqQ9Y6YQ0atFmiZn+Y0QQUHYIj0Fkypv1DvDFOjVY7BLef6Tr4AUT3xSViseWAJfn
cprahS/WXXngVhcx/BR9jdO6gXDsaVfBzF/K75I2NZjlyN9QZsupVyaHyumLZeWLmpUal75T6ZfN
nEMWkumLwDCfyqIwpxJMg2fjTxug8b61priz0FDiLWuO+LuO7MtljeBxjaE8w6wwDdvkOmbFKeDb
P5C446+a4jPDaEyqNR9XPCcX9xIs8WcCMAH3yNW8kFiviAR3aXxGCMRyvkkQjw32fPDXOuaUsLuJ
ZSM3FJPC43Dfttgqy55NOD++P1uS/75I7+xHEAXeYDOO/Ia1qENK5atcuj/RZfjO63rjQmpUn24F
FlYToVMbaq2p1BxMwjHsVa4f/8Q5L7I9UXUne7NsbZRkt7JlVeqEgsSOwCHo5Cp4oAXT9zxmjnFG
iJu1TcRHiOa2dSs1KOz5KmDJxxC0GMyarshhqGclsb5qEz/btPLhmPxHL0L9ESFTyl2xaP65Yk6G
cZz2t8dfLOsQr1ohu61Pqj9Fq/DyPm/7gk5X0+8v+kKPC7BW0+wPKfBc4qzO2ZAWbsvjtBwVHuFm
OYUmQIfXEaCiROo716/51QqnHEQnKuIzufpmCoEFAzVmCMOe3mmSdlz2kr+3CCnLdyljJUwRCiE5
FEVlEcwcZ0LaegTxT4xhlhyNj+oEqrDc9EWLTX27ZKZCXvvW1XEw43Fo/UFXCVP4XK+vmE4INt26
vtFaEP0I4aRoCdBXWlsqwLnrLv0A4BNwRF/brEMU4r4ZKqkpYjMTfUyy3NytUt3aVLVkauP6BtG7
dAg4Ebx9XzoiVYV4s2j4ODQ0oKxMZN/wgLfNKLUqBqltbscTZt+NYgn3hTcBG+1pT8WUTOaW4yA1
RIOSEGyOyIW0uTJ+0FAfppOL+IcqRZC/Rxn1kV+THxZTO6Ofmn72jSn5yLLojX6m6Bi1hu5GaZEg
at8aTi7TM8J15+Exa2KOnaZLuQDkzA+MrPdZ4VYZ+hPvH8WoA5GV7oiUYDVMcKwhjfruWrxYB4bS
5m1p1y1CTXrjRsyM+rKOSV9prn1ttMGnMACsbzLKVEiSUErjeNreOsUhb8DmWc/dNcPjACGnz2kJ
y2AltHddeDB+BQJMrQzaRLhLpdMqmfZ7xfisjcXtmQR52Gws+sF8vWdWNoBO5eDS0iQHj8qnn024
e0fsp1wClacEt/qWHPTZK1k6Ac/D+4r7FZNriziKhDDL9vO4IkvxxnMdp14zpvf6yhAt4Rxq9XVq
ZXCkdCVgxtd8koP+qkNlKECV2IYobrnwCqsuRwH/3yZlRDSQebwV/1Hg05LZAqA4rNGn5NTqHj39
Z4fDjdXFoyttwM5NYAlvjwwRsMIf3zWlhr+kq1wQ7efLki6Xyf6uNEFRgDAUSMjW6SAu98J5sJFY
jW3BnlEnjXUMBucxPxJDf+jkvnI9aJzm+wwo62tFAjcVF9m768uAIWAdPZZkExo3cgg1XIqfZftr
cCJ4ckm+Y0ikTV2q124Jc0iNZDSA6n3/YE9rmYwkTlLpIgTWDex+LOwMedEjj3Ewm4kXIyDF/LSa
qOcW0SeauhMcyjMMIHczgsPSdN144b1uIii7/0VRsYPtJBZaQ5c0G506WqcOVfsJElGGa/dkmiX+
F7wshCjv5gOMBOoVV1WdqGyLcD8ueh72m88tG5W89lpq+gPJOoS3RmfZRZvYVm5xD10DDLEVi8Mx
HpEtHi/BM+T6x4zkjTYhU7W+IC4qYJSe1VDu1WVod7iHYfO2jLGYrDzoYS+jSdZywzTRjmu3gm+h
dFZ1bpxq/Nh21IB8yqBfPBvfSKdNxEU+7hLWsihy12FncahzcZlrIFIW/cLnuMCecykRPDAK3CYi
geTWN8rT061VfTcSFR0epFNmPtg+RRwNvTSgzsu0u/CGqyJbjakGqxNmacm7PVMvkrtC0w2U7Rzr
meYU/JRdSYjnItzgy1DeukhAOeg9SsXMhdZ0Mbshu3J7RZjUAQUIqOCIS+7hp1Liztw/k3ZiWvtk
9TP2d7OzjqlZY3/2ZkTXKN9JIgU+DnQqHrF4+snif3/4Z9O1MfS93+ahuuTsOiRXeQLxDOcXZRts
vNIvpk8B0j1gqIb7QR7/gfei2uisA5zJFSJhsA2LzTWgUslsAdoGUnBCviklVhm9+Pzq/wIJUfSo
FyzJQ8iqiBMQ6DBKdlYjk8KJauuul3ZVxQ//p9UraYcFpFm6HFvXYb6YGnrYLWV6nVm5abb9PSZS
76jGSkOkULzbphCSTDXWWFGOpDRWMG/clo/XQu1jRICpZWIolPBhC1jRQA1mAE7b86zxRIyrOTWs
OJNgaN1LpZmEd3gcnTLzb0d/FB3QsDXSQeniWFKm6m+JOY+EeBHsRyZzQ2aitrPsztuAmhgc6/3o
+5d31nJPEYBNI0rPd9qAv/X+vtcozbZy/ONOMWOHkqnFhKLGPmJ+r3arqrt7poih8qcHrvamVPxi
TQpb3o4UzUQIum7lyb3AB0jDDpXViHvtsuhrk4vt8tMMw9IfoPc9SU0PSarjjNv/PDBUHOFFTgVw
Rz9DjR+XfRjP7X36tIWjaheoTmDHkt8vLca4iN5AwxBpik8pmzfKfe+Ng4K6GytN4IqBWIITU402
6hEp5OkMmChaDQJ4+73WzrcQGAdIWHPxddcVdPJ7EiJZLBBiDLoaJRccPAIbio00Chr7P0pJ39+Z
GCLWd38RjSOqPukpDLRJ7gcBSNLIQwkGPPXmED7RyzjfGLtRu2s8nY8g2I41EonIM8Ku5aJLYFpz
V9vEn6KUNRah4uCMrCnDQGbHesg4kx+nligwuBMJ2Z8689710ebvr7Wrsf+Lhd1qnd6MR3btmalR
UMeSZcdIiDM5y3SjZeHJqZS5KnD5G/X5NDP3AJy5ITTak2w7KuTZIOdQbzJQekPJR5G8fh06Lic1
v9QZFfZBbydwfN84Hg+8LWrbrnJAZ6nKVRyVqg9aSGLGBk70nFvJAqfttDUaq2jhESes6JolMGx1
qY+rcZhc/ZjMGhivjNUlmv0XCCr9Pe7qz41kYewk/OI36BwXthjj9SISxTb5XvpNNG8MfkXeUpLU
8gcYStVmQZhv6FqgizPpj+uRpmnN6JNV6gINjMODGlJBDoeMunDR4tagBIIShYYclq14TOkdm6ZS
SRcJeQM/PUOK97ipqeFT+uE5Xl90Z45t5RSZcm+QdwB6bRZRr2Ia26WFFAh0grmsK0xrhDtv/9tv
HP4l3bgwQf0iTFzbPYTVLUPAhhW43Lhoew97wx0E/d0N6C9dfk6dGy+3gYguThLtv+WZxlkhtOg7
AOp34tr7YUnkVQ4BXPw8IoqxKHuv+AoSyNg/4Nz1cKsuTAtHs3YDaI3p8PCGrsvuRUGcwHv+caP7
p8S7lZJDR1VatIGRPFz/JPZRlplakabEXScOI201oc6bw4475n0USQZosDXS4/9s944pScC3w1KW
N4uCB8Fn38qH3lTKmjcgGjD+PgbNspgVTAvBEV/4EyHXPa275mDY8Ww6B2AB6d9ARYw7YX2JwNPO
M8pvz/fwOonp+D6+64vauJo0azhKUBJby5yEDTH2sar6Uiw+ggmScJrbONNdF4DTLIasSQ1gl4iy
knGyY9yCllhw9lGs2C0hJeILD0FMeOJSslNqeEO9VaNarip56r3GK5MG6Aq4F4O0wCNlpSBOfDs7
/RWIEur6aZPs+9aXsxICnKAJvV131h2BCwAbth13/S66CTY8R4hoK6Ps1kgESVUMXEML7Xhu3Kxd
tzs+qsJ8Sg1gvMqwGPQLWDMjoZBcbTmLbjOO0tXttySwaYZzWhxKt2u1HqaZnexFtSGL4veaRiTq
B6NdwC78e8ZYSaTPYKMcx3rOh47RDt2l5bD3rmrz0TtlSEHLowI/JtXQilQbZiiJ/4ISUv0O/qq1
7kIjWHKRgdh13cvBSeQ4Ws3/i0ZNbwXoGzkDUg6j9cOVvtAA9USklOXygEmHp8IEC0CrwKaTUTPZ
QwcGoDrilImzJsQTUbPkCarQ+MNAvH95mLgibCHeaGwwD0x9Q7C2kzNnxV9QNAqrQwUJAOCcZxhS
gb8JDnUMh9SjokFCBYfuOdRxopABN2kOQurYY0JTKxL6oM/BYnsyJUAtSjH/kHmhS8/Wb5ojFZEb
V5yvwjsfJB8djpQsk/SVX/BhnQBUl4mB0YRH1Hmfs1wpniaivY6eIS2jP50Gva9BONbPA4YqAmHc
3AM4+QzN9ZijfKe5QYN3vlVPMWVbQuxe+bTc3HXnbOyYU9aqvBpS72PQs3OwgZ17OLpc9MjCpQrj
HckJoIgYfyye3OyagiV1vwvrqiv5uI5+COf/JXGo0AVvuVdthAslnQEeHyxO8UewFe5tMOjECGWe
WOmuRVj5u+xn3AZ+e1uIQ1yzVVGzYpe1jNjA6R8oMZHGptwpyMg3I5owNrDHb30q33X83amchrFQ
XGTTzhl8B0O3qHkkckcHhnWMjv8vvCefX5xTNlIHbGeLj3w2S77JZlvQsoqFTj0WY5tueTqIHn6G
3HWdz629tDcgZzJKjadb+aPEICu4esigPFMAtrR6xnjirz0sDqZrFCfFbBOog8B55boZo05uLXKD
8b8BUlnAtT4+kuESOteFQ0oHa46Bb/uOBPeNFblFjpgoVG0ERPuBEITwmo9KebfYTYeINH0ortah
vI/m1f1VUHAMOd39RYDFPD9Gc6KUqDldrUlCrQ3cTQvcTn8FYPszZygTmtwpKOpMkmi2xBOHhKfv
qAyvxwmxZl/bCszdikdukL5sltt16gwi1dgyCGyaVSTPqDzk5oLa/ckOBm1n6xWAJJinVXdtBecA
Bp/dPtxKriAUwXw+OfJQX8E9w8R87wyguGoNeM+hLcAuJFirYLsgwcdf6RlWjyeMXCWzftAI4TBl
V+Py/tlOXSLkw5gbpqAvIriSbBFTd+HaiTtekBVWzseKRvJIYsLOzUIii5rvtEGX34LPTczkWfZR
PvSp/P4jAs205zagKuBSEnGWwheVaVR3hWsMao7fwKUly96CWlnrgODmB7tBI/rOWy1IxnyawpVZ
x+ayv+1f8DhHN2ZecHliOq5CX1S8nvBV20l3ipGCisqGWnJc5/giNjQA0hYaQzGFm+eK0SPEnCj3
uDkS61nFZl+kQq0YQeXMq6GoFZvh2d5lACkEK75iv5ASLvmUXaxfM2rk3ix4cseD8+rf3YTu9qMv
14U5MFxbfIz6P8tSBlELR0+pcBnJsdrcpdDN7cF24aPFmGN8d0gsLJ6rLgP0BwSPGwg/P84IiUfv
ZVvL36004mDvmT3uP3UKKXBm81J2UBgiE0GMmND18zsDKsaOt1O7KjbJAiWe8/khf9ikQpeoJxvD
Am+MrdLN/OkMnPp8oD7MMKfRtvVb1YayrcHnUAvoJBVmBrgD2pv8SOZAWKDFqK7jUQGEcim734mK
/BRAamR+An4wVjbSAZUeQNP5lLk66tmP+cLteYXoDd1EXaPicTOX5VlAWthNXrcR7ntZR/uSVd3y
dlWJwDaR1SFodHT8L5X/lJt+GFXEeT99us8nrH+ccvf6j6KBdUW/ekQEEk1b6SrQgqasriOcT3bV
UQluQy00ymKDuTv3zfVA/consu2VkTYbVD8xv5phbwdxr+RgQdzdXaLms9UlpvuG/5T4s6kL5Ord
maGO8d9Wa8ExUwYfIKpjU0V6YahZ+TIVMFH+IDWLBsgLCKXL7qiwHHStXr/CjggkV+a7RwqRFs7Q
RKfIMNRCVRndgQjYldQqFOnsPVkoRnFW/XN1sZnGz/8/W4Wxvyt9ShR34X15+Ca/VmsxvjwfmxFa
uZAOBP5neqxSkMv0jPFuIrH9eQJPgmWdOd5vxneWa6A7JBODb8boJBOHMjIGwkTwP3so/K8kZOas
NGaGdVFXd+fFyRz38V8bNqwyRTpJVX12fU4yXhAlQ0dp+nLoqHwKVYAlZ0o4Mw/5wpmVNOR7fOf+
lO/Gjr8+MQZp35QLY2+KZBUHr7YjBGchOepgoqfjhGgPACJBXxqL5nSasASefXrFQ4p1i15pAQu7
A4BDCanM6Z3ycFmu/I9IWsijnLAnYHawR7BMQYAfric+Yrj7MnEmrnmrhU9tVwp/zu/i7nevzLJN
sdLexYSOYoPMTsrDSu1A15LhXqIJduwaabSoX3WW9vS0tYPYBlC0jaxQA12Fmj7TCcg4TyQZyQAD
RGugDx3zdD1qJcPtFtEzyNlO2trJ6EiBdtBIAVmXPmXGTtz2cFUhHsuLuq11tt22CyQBhcXyxJ8k
5A7SvUF1w0cQ/fcrv2Ak6v76NOxXKDBOsANsStlzLYZRCS/K/Zl1wdAMeeKexlcLZNwOLfWPoPI4
9BLhKheOkDtSq9BvUzMvhmDR/0LAa4eJ8x2Sn6+fE4dlOK/Y81fr3IU1LirAYyxU897qp0juB0Sp
OBED8H+8Urj+rZAQAFmFCcWCcGjmsE1LNzwwTmYUBEpuIC1rQJCAIHG1egP/IjhvlM3UjncgexYD
ysWKDeNDOryoAtsI06bG2lI9prwSahiXlA9bHb2WFOdA3z4hl00C930cg1p3aX2xQXx2PUyDXfmb
OlNgOxfae5U+Rvg2iDtDzdQo46DoPld0L0+dwMdNiSKVPwPThBoJn1QrUxyOf3INh5DCrX/D1iHr
25ifcSFEjhlObDFi7oaFEQjIjOSvN+cavfk/J30a3yFHA3HjUQnLlLNKgCNOdPeX3d3+F+/QOt0G
CTx3wcYQcke61J0TiqNiCTQ5npEPLdm0Ei2GnSyyvepb7/9XeL+S74uoecoMDyRQI/mlfUrjrvIk
HocHxJNzd7cVhl19AanPy3Zj7qahJaHYqtjnWGSdx2I7CCvat3sN/4GVvCjKBgHYABmU5Babghmn
LlCjwl2LCUmMCIkdP+ht+eKrXcXvneGAqg94eMJAMAgsZc4TrNit8UKSrm6Utn5EorjjbF9ZG2LK
qIWIf9WPuqJ9weigOwOwiK6h5NsMo1QzPbvqGZ6y/indAqS7pJmRJ3Fvoi250b3wd4GfGWU8HMCZ
DUdX7TBNnTj2BEYZTu/F6MB8Qv7PGyAN/L/snMfAHumKOR7zUerrIvlSCqo412iZetE23xUF4s8z
/DgbDXIVfXCWpfOp+ECb0Hk8h26WRtTvpg3zcv9wkZhktvzrReNh5I73Bng74RIa62RtVHlT1j3Z
soF2FQhMz7hs1famkjZje+6oVO1O9ITdXlF4W2RrBLQ9RozBs0SvDoM2W3LumZa0ordJR8fQ1pAh
Eo6lfKe3DCu+0mdzHgC7cQL8gpJgC6RgbCRwdl0UnfjvV7Ze3M5qqIZU4hiCN1gVeKsZtzIIVn+z
K2akyqvmoulIYrvm2G6dgWKQ70sg5DMYIeUjaBke7TaEM42uMXCJcQQlSukUJ6DXstfMUa8IJ5Lh
eQtfvoUIxbl/pd2d9lBh/XRpNhJmGJLSs2IlSZfgsTj3NAxAm1Asjc3/6TC0YnxSkQ0jlsS6Bhj2
WYHUBnl9+YUV91fzZu9Whwbe0PBAwv/ehSdqm/7NWkeB3zdsM3vUBlDG16j6mf5xBCeFXBj2wtWc
uXd5yu3FFjd5kEllBAOBdat1YXMeL4A3SoKUJXMcXfyBCn2rXSIW6pwlBXtIqmiIHbCzCW6fmPwp
zFw6jy/QejlYtbbRzg52HcOshoHhZjfKYrkCR5PbW7zVJRBmSSZ6JtVMsePCy3hJrDAoKbF/nhfC
dKTIaC8YdpsyyMGydOLGp7wuPwA9X0NOIXwDdWz8InZjmjLSy6nyjqyjmwS375Kui6KUf4LNMXce
P64DI9I3LzTZEV0i2eglC21h/eyOmG9MwV4jX83e7rmMCHS4SXlTH3Fx+rliB88iju611vEHPhLZ
q9TQ2dwSziiIayPGSKAxEV+46RgCIF9lFMLkiIGqHLCuvRmhs5sUad/zFGFNwYkjzXARgzPTQnrl
8gVe1tW6XwSXFipXWhdhkH0JCl05NkZwBFVzxYTSvQLc7yh2qfN28aB5KzUcjiajTP2tA7D0oKAV
v4zEWRwYd0W6ZuMIecCyMIob17ckAtrqZqBUiGOZpxAl6JUCDyUc1lbPZwzPY6V31DjwCLroYD6Q
OVcIQBC6En3ZSsSCCf3tQedidpS6ASed4ulzWeohcu+IyimIEYBd/VRZA0txQ8r3UxWuEnYInq4V
quEe8dmKpv6yTDgrqaRiNENGVBe5p2yFysz4EfP2py2yUJhF91/z5S3qVCiWXFEdqejR75rJNTIk
tiOeREUtbk2XF+g4ztlap93QLRmVkXsRdgKyowbrVc/k00QFaf9uJKrq8sPAL5f5FAWjvwsWkGHn
uvbVkRFQzwAAypkLIFx6OJlLGUU5nxPmp1UWtf+evmSd5rqDfFg3Nx5NXVBQ2iTmeqMZk5B1du1q
qTqZtCRhRUk2+WF0d3zjWbZv7Hx05hWTsoNIQicVWhATdWRHXdHl1XIwR21ea9/82ebJ8FmNrsk5
bM8XS4KzXd/QP3EoftfAPpL1NK+t00xfWaz0wVzgHxxW396sIXIobxX0COj76DzD/mLp3+3uAnwc
aQtWKn5XY6EOVFyrAtj4reW1BNi9oYK9J5j8/KBXpQCjVoO/aGKssFYig5X/Ymn4Q2WvBvrHPwvB
uNTVFQnv1IRge9Mi/5mZrluxqkKw+iFXOz7lbUWGrUXWVZ/l5nHd4nIdfV7LqV8gZNzTdneeIIM7
YEB+OiJc6MEM3J/puw54mRNONDzfx11H4Epl1V8b5GOoSHjUu93h9yWNWAlcTwyXN+HQHVaw++zf
7uDkktR3xfZhQ0D6Vg6g0XWtZpUne4rS/+v0JtuK47vJ3HXRY4dJ9ZY1a7dNDdK0SgFsQnoi+DE9
Px1bhgxcIy6khk39dP/CRA6z6qSFCb/8iZxqDXhF4OIO7ZjEqy9skGKkMMtV45r6ae1HLICBryKj
J3QlCQr5bYWIYZ1x8Y9nR3EJ8mL+/2thvXoBZYDS2nnkO4izuBm5P2r0li5L1G00IF0VpBD20gCy
Cxk4M9QS14JhSSbXJSf9auPj+btW6t7scWnoMbe5XyxAgrvjnUjPCJFtmpXOeDTeHeZ/i4TJaFr/
tOtOpxEuOWiIzfhpm52BwdeSCgOpBzarUCcdy9Qvs0W+3cLoXS2/LY8QtxZJHgPfmH6TgMu4a7ch
8LygWF2W5mIAT2ngI+jpNK8dSljtnHD6KMD6fUSkmGe0EyAVv0Y8Uf93XIMPCtJSxKhuV6RPB84M
UgpaDuGa6Yu9F9MhVD+8G8mHah43/FjjAEi0gw0zUkLqRpnOm7i228DlsY8Q3dfrgIeCjLFftO75
yk/NLQEOJnIz8S8lj2ip0ULNW/05VUArHyjiH8iHvbp8yXkZBe3wHVTwRm6kocph8p1BC1lOM0tB
fTHKToGF2KkuXCL5i7HLxm4y17AFtMZuw7qD8jLJWRlRYu/Ub1tKGUyUbuB+zZivlhE6TFdWOKBn
ATqs4cDLu8wHguQJu8cyIhAZz+ZMsuJEolm6T4avG2TzCXd7vPuybzGKWIE1Z0hlQzEfJy5yVKzT
iDrziY0AbGzYeMAsEc6B34Q/BgudLvBnTIvWDRMe3I0kxyGqppddqlTZMfG7rm+aePC3tFb/gSIY
3TYIkxAzR18qXoRu3iG69X9BGnWp/awOPON6Ho2qGXT8UI0QFm16O4eSsu1EKVpfRf+EWVQd2FWt
Omy6ndLSprXwn+/h4yJsWcj02/v994VAQDZVWwCcEKnmQWEQyZ71tOfwedpRqpWaCtFiq/gJCKzP
GpP9BbmleU+0J1WC3tT/HwtA3vAhDmc5ALGcjN0TAp7dpa2Bj1zXX4AJB7d+Fv+AezKNX5rTH8ac
7KuZRu3lkNuKWnnz8T3//9YwPer7VksQ0nQ/YXd190koRQSSD9vffeV2FMi16dvE9bs3xjazvth7
YyODtnPM465ds4Nn38GPQggTI57ziZ8RfCS9rRJuy665VXySLU8k4+WFlGwbE1N29B+YTnB2ZFWA
f8yLiHDjnDxsFqcW8HWmQwy+/39kT6nJ6kes6cxYa6bbMvccnf1AEdsYvPwLCivTO84zRpTL481f
/MoWwi+5ohJ3+ZP2xWMQOkvDqnw6AKthG97nHtmQgFv+lOb09bYhDc2H0Uw0duFjKmgVEhsKL6MF
Y2vYF04gbR6WX/+K5YTZV0vK9/QmZfrjfAH2Rhl8T2fdZEU2Libbs4BQvuybyU3MUI4meAVVQY3E
qcBiNBXS1zik3aE2J0ZNaBFgjsJRk1QFmFYep8eaplBaeABKWQj3PsDiu8WiFIf4TltFwOfyaNpI
tKssLQiyqox2UjQmF/hWRbJGYnph6YxC+65sMYdLa8WKcv/uOBgOx6dXnfJEa7uv7QsLJVIc/OGV
pXMwqZwYHmScrLIZfBP1/k+IslePBVgb+Nk5lg+rcdu1Dl9XEOp2H0Boj18Ubq0E8Et7RIm0tfgs
UXDP4fxwc+LkqTXqMx+kxw1dnOpkcES+E82hP08e/VbxlUVnfMZp3idklZAbyMcvl2wo0YU3JC9s
Phj6hrEwamW9cdy3gPpBBwfqRYFl8ZAwWYYUPWAUA1jubHyQqtNMrirohrTuZ+MLcPQTvmBeO6zp
f1BETk66PIckEGWiJeI+cz4xnP0cNUCo/YrIrr1/YN5aCJsOOLOLboo9RaTDaNB5VZphRTRjHQS/
pY24vNqy+NKtgr9V1jL3ZJ+ITffdpnotYk8QtuKOelsjkNvAceilwez2J0EC0lUQ0r+uhLdXYpb/
vjihA73CMTim0DFsKvzDmZs+h9Q0slVIfR4BnSbJBz2nSE+Z26n+NhN5zxLtM0kUb4J6uPHOz5WB
VhCLhyFaRYLZdUnHBazvty5JOouDUgtOANJ3OBJ9z0ZYbdPqXI8zn1s7A2bnDmxCjjyIjKZEYulB
FzkUJI4KZaKqi9Oaz6iIg1UPjOA6y66SxQ/uYCwSrKHV781UsyCJUSbCS51d1FxKGuTScqNIIXEp
iMZWb7LzoU7H1gIWknrsaXjc24Glpgr3fWEWGmCTtypujFEQAtEQmZQaW1Pv6tPokaA1UeU8Bs6M
mm81Ie5ZX4zS3OE9EK4Qi2Mv0B0m8Ufu7ooP0jA4zTZOt/W83XdLD/IkrIfGlW6QsRPKJrpPIF6V
fojNgSXObMZ3q13l3fi/2KZ+ZzIULaQV3RQqCqdbcXk6zkOxrO6Zl6Zot0141jsp9meIc6q7u5so
JWF4+5IQGr/6bx/tPXrI6R0xVVsMX8XCHUjwCT9NZJ1vvPKcEvQi0beSt45eCRyn8Tn5DltQadUW
8BzjwK4ZTStTl6dz3wnipMgmGwF+COrSbbprrmPewoUqWgAiGjNt/4wufwJMRPqk8JJBhfskW6iC
KI2Qf17f0stEnA+zJSs2m+Hi4NBcNHqNZgpw1x7FWKr/ZfQ1VDbPPINwlRhp6Lkw5crTHDd7+uGd
31D3S2IIf+XbiwaDYEHoh4T3QLpB+31mVs5ZbgMjCU2gxkPCTfRc/eaHNXnm2AfS6DcdenjY+N4z
u5dDc6jt6cEUwLQI7k0Rf6Xn/l4pBWBTgun1maggVCFC1hJF/CZeKm6JWAin27wjf4urdTojh5WG
p/f8VnQwtGlwdKVII+SuidfVw4wg+iFM9gsq0IsLYa5rtA/bJat7EiExtw8bwtxxerQ4EKKlzAvi
Ym/Vi7bh3TAstiGExSpF19yz3dYgSHqENvOupTbg7rUn7w6EByst1lRhLANp42eVo7LUoSIVBzEO
wg79N1VUDy7Mv7XDvC9wjarV3kWoFUXd67fL2lFcKVDCDgYye5gW/rUK6iQx1fbcSGLqpyT9pbkk
7Ai+lr97ldjH2drRd/YONEVrkWaqWojOwl10zrDnCJ9gBE7nbsTeoNJf9LxFen/5HtQ05fWKYlyD
MskiGAg1h2ZavAwXonDtgNm7z+cjoyegqbjDzkidNagdDqi/b9CTRJWeMql62AxlH3cgBmYuVAdH
LG5CXyYyzN95/xU70wuHouqUG1tnhnCoBhuLggq8AbJa81cheoBMpow90vHbd/ASs64B8Df2mQt7
JgfCgFPzVIcwqzopA5spvLv6LOOiqo/INhzL64PFGQpVhSEGkEP+nwCIIYaphP0xujLWxMrfHZ8D
oLyvTkbouevzByz1p0kYh41fJnyNMPXtnhOSF4aXlRMl7JDBcMQAuV3r5s90kzBjDOoxpaf1PQut
EhaVSu5LoKyrir/mSiijDdyyQK26U3Lq3iFlewNfBrveQnHSuROEou9xqyDYbkmO35T2AsbydSH/
pPuy1+5JMWwFMKt//WTHjxHKfCQm2k/UH9nG2ZBy7ZP08qoLV2bHYNd9NKscdqfqB1iMaahpa9V9
GS5uisWH6LOE95QJjVnB33M7YYg/rcTXFz+5/8wLQPOv4uh+gZpHS4JnWtPm5R8Rhhx7Fkfx4zW4
s6km8fGcbCHk+pBQG0keXLg3wMCeOZFyIQpHVL5bZnYoMd5SBaldjbrJG+4nZceAV+/+abHu1hqj
oajuSSX9eL4tktQH2co5gSoAr6jXSr5r2m96E41QpQTlgvG8V+IlQ7/ZC8NLNF8zX+BBlm044R9F
S1GNtjghszrFxty/DqmSMaEDzoZ1MehbUXDGk7i7vEq1hDCfYv7vJH/3BIdsOWSNQtEv6FXDZ5B4
7wd4KXRi6Dv8s+xAabn3zFRQ4I32PHMl1DSVNm7mFEYIQl1RROKlDcJgWBKuHWoqAqbaI+hsOXoR
ezlgPSned1oazRNDywE+2gEn+ogbB2v4QIVzBrSuCV1dAIzBDS+Js/HH8ffNiluNWDNNXMQc11KQ
Zre2FsnphhmmHAp1VXpNP/X6zER70/4R7Ze30OS7pUtGxQQn9xVSulCZceitcDocFXWvINT6owGd
ob9a0YK4YFUvGdcRAhtp01FzT0nYZxChc77ksAkwXjbY47OXLgbYV4Iq0Lvc46LLdgJ6mGljOXeL
z+RPVFSe/zQMHGVUngj1r8jdS1f9OAI3kIPf/ujECiIPF0jMYqXFpBGH+e9cmgpLk8GSQWMjM6Si
vptfHMNKLsNZU1kLLSJTT68Psf8vaPylDRGNHqkKEHPXWZuudP1xmOyvJnX176n7LvAztsd3kkKt
HcXy9zI6dEPAxnq+oI6eFsiOmr3W7WzJJUrSRz8PfG072D1hsUtxJJ5NzjDKvo307/pMRPqTt61r
TJV/LjJIqfWJGKrbwkod7664/gOk02W6h3rl/lVDfJyGvO7PX0qiHnfb3SKHTWyIgp5eSOjhEZ6U
RTwwoJS6ZEU7q+0a3My7PwHv+uHLxC02AMKZq50W1T/xg5B7pdewLhZq8b4Ll8Lk4dz69ALWGsx5
pLJyMsX5uLWKcTj3wiSDpVkRFOGAUxMFi/NLNfe6ym0r6Zm1iuiZXMODSnInS6VOp0f93qM021Qk
HBelOBQHlnM9OEla9e2kYdDRAhx1w4pgqiC/l8VDwkrkvc4hGKzJkH3Bu7+bkbvmJ1G362uDpUmZ
F+5y5gW/TFq2D16DY+SYI8eR1x7UXuKqK2fSub4ZDhJNlBNoxwJjqpVZeJUhocDOkA93PiINSZlt
8u/BRbk2HCUCgBi0U2gW4ybPPa6pRIMdCmlqLgqW0It2XI+Vn1Vb4PvfU2XcFmxvm87QSY+vM1Sc
bfukKBUCbQpikOKl03qXO7noQ8xVa+Cb752OOJs99Ml106Yt7HpTkcgS7kxz5oDaM1yadGbLsePO
PEOZ6fYaXxD4paZDWVVYld7Ea0a9RujzXJYBgbICNZmfmsqW6yEOGAGPaRp3P80i/KmkHrqPaJQx
eZllxq3afPPKKP44N7DeMbj/unAphzlkfh2qCn353bhHZxzeEjbd44pkoKLIbHlmd3F/bk8Gewv0
9YtpWC6HBEikyWJLXTGv645SORGU5JiYKh9fcexWD0A1fAFQZv7pSkSt0IXs8avMYJKOuzRRMHOR
CQCwDHOI3AvL0TOzPZvK6hvWemHIpL3kmiTMMCgQRc/l+6dZYbejIlzww9gbT9aAL0MWrvWz65Fu
gmpe1l1RQPHm9Uj6UBffe5mhdW8Kgps7rvhIuMWq4Z78DQf36yhpoHKwAKYuMFSSu3Xt/K7ail7E
/VY/Z1j3zJ7bIh0xTEDPUbVWvklxEqurPaWUcjImRkc/1xC+JN4YsI70BbWGuP9RUFOus6r6oXTq
9a85/bnQyNG3qiq5wnY4Qjp6gdalJD/WXyMvitR7Vmd3bziVTUba8S6XzaUEYUS8n8TON9bApOKI
f9foaAOhSW+7X0+WjKA/Ll9Z1jZH4Z0MctPYaeemXm8FCJlKFQDvtBkh+iYHAqRFqb0jutsGiLqC
q2TIJ6OdPYxIipOi45fq4bYzht4MQb7HUgzsx/uhIbUWDiNg4RjVTTqcfoH7vhAoMbPDoLDtDN6/
a6ChYH+Guw01zPbu1sxN3dllMmBGq8/LxOHg/yqcY2CL7ccHGGMpxY4hBDbe6T9LoKU+aLF7BORT
HF1yG7FZtrHrTOL/xSf1y2KZ6XpoqinM7p+E8v6MsITgIMF51OR17zJN5/Z1Nu2lfr7VjN6cRIg7
Y+wfKKScLspy2ujsbWM7W1eHTsI4/rQwswkAncw40JKdJqmDr0L7x3bheny53Ab4rNV3/+IUY2W/
Zxk/cxESzD//YNfLpxwvqfX6b0GMKQQXqi+lLALPqLyJHqp89TviMRo5mauL70S3P1d/MzOROL/p
51osoM6yttPt/pXOnKzU0I+j87qleUBhm1vhJKP7C4aVYIN9ynaVHHuAhmqJgLCQCaGNfhpgm6kS
5CpKCQ3TuD5oDTBnA7/1dV4euqLhdqysk56IsKuYTDt1khZsYsijOey5oTRfUrvD1FBYRr9dwWXS
iJfs3/e1ncbf8vcDBfLGsaPkHo7zMKPIwUzu1bRurDzDcGtRAq67W0zBMLu4D81+6GHPXHBTrXPB
AlaaohCw9mXjib9SQdDNuZNjSNmch0XH85HuiEz7bsmOumm69JEQ2CgfkQjzB7VM6eI25JzwY7+L
JHhevRdNpNezM/Rxf3Y2jQp65XKl9E6xOt1M5uqS7TXiJVHoYEVF6mZwX2gAIw9Ja6qgfRm+zi2m
Aelm4k6i98+y73Gf5QMP6mjKNuEkMl7O3J7cQR105KVDbtCRjiOy5KS049oHCWcyXjFs4vGExfTZ
Oum6Qzv+RJVLCDqhAdPOGDB9M5NMz5o5fQvDMVkPuKnlpbnTxqHL3otB9t+tw46V/beL8AenWXKM
0qUzbQoTkq661pjE7Y24TVByrRuWfGScV70esVu3bJBspqJAocU1XUEfj9Nsb9P3Q0JLT1t9rWaT
AcZ7d7imaa5iWpTnJ5IpxzEthwcF/PqZxxiyS6wBOzahB3ViuEbSWmK8FUwVktbV0mxQs8geAf+C
blqz8XMB9Rruj+8fs+stx4SEIy9Nrg6vFax2KCIln1Wa0ROU4Fz/vOAVc634wtrkTcHvW1yHdWid
A08QyEeCDcrIfSvT20j0ix4H4LTBhGvimvxlP2PUpJguKGFjmWzFJ9B32l9Va/Ag2szNPZfR2OoY
V2bkcnorKzUvIm0dwU20xDCitE5EyCvBWd8PN5aRwfrBMymohEVLIZs6eDOiXzrp7wKOca6wdkCp
shNnvjlqsFktoEAL3erPZ4Ayzj9z2UHDLs4ivS89sLZl6F8+JI9Z0nCjf7Y3jEijz0WiBsyY6F5I
DfcsVNRCR/JlQIJGr5V+OvYFKAR8PcVlxGBemgN45fSSzgMAqo4j2D6PVfXpzLmMkdp3BBqGMPkJ
JWmRh+s1CvDaUba5IDp0mnie4nj/UmXNpKCSoYQEvunuslkVhuHz27QQla5Q8pvAD8LuQFJbb4o8
VR3QJB/0oO+bQS3pJzHXL61hGAJvD3arBT5B3HlbOxAhn9MCgGemrXUE5P5PDS6MqmxHslg2Agfb
8wlRi+SJIYhLjnO8CEmfGYe0emnEK8WkcwZeEiwIMB43Du8qLii7gJxa6bcwblxb4XtyWYOjRdLi
2xIlcN6TEN0pSxAzXAWaOwoO35ZKQ47mDiKHzSLufvxMMCL0+49nw7giL5+WhJcsvRsNJJaHtmjj
ZKYZosNzzKdBqvLwerFZJRd+/GgflvYgHJh9y+b6GEs+rgI5xl+21HOU4tCwKIX2BoZKrsk8EOOe
ah/ZzX4JkSstUIeNYnRWd+T6euBTqZqXI/0e5ZOesWaQNT2WD3sUgEaNmdzBFNCNmeYGcVU+Yeam
mpWZ8WI22UVX6wDJah+XWJ3Dg/xUpLZRHP0MNjsJGi7zGQzA9vubjJ3wmKcxThIWpy1lt9beO81Z
GdFEvFV1tCqcMAR8GCQnPBKw/CctDnANdWlNVrczxQxwS5Ahmo49ePcmifjmJsFXXvsCNS9+Og9z
21TApMvBUCLIWH98Eii0yGEWnANYj0Y56dKWlS8g+pk2UXZJBlwb0PXd5Bce2laHl6B8hih5C2/b
FlC7AdKt6jnvuJO+nOs/fT2fGCUzZymW2SOOfPFMR1iD+LvspFZvhB3AvieHOXi3yF9etNiJwHbA
8veesfYZCI1UiuH/ggzimm55JKJ4Uy2fJEhNj7WMwx/O7YYkDGk2YocGEUSQZ9mIPM94RjNsgmef
i1YwzWT0ySAJG2bmv8qtKIjnJJ7iSe9seDc54lTLlllnmtgB6DVWIUGeeTAtPnJ/WEFnXdTGh8SW
SBmnL6sTlfSvCBScIREvQsWa55Kv/3d7BDyOG2L49ll/50rkCciATqxRXFd4T66Vnaa5gsYMJ9Nz
EYzBsXqul+F1omHo2+n8eVMur07kHd4qh7qNoXTwAt8mppu7n3fPG7E6L8UXc2dx1KWLqXRSnLiS
GN1b1J+8QbZYdMGLKsj10EW2IBKKfw8XLN38OAGPSa6i/KghNycSByih2oZhh62+C8PgmULjuNUx
PwVlwyiwgpAwc+SVrCuNgpscJl26hvzw2iyghFyrzjqkfADxB7w+GhaTfGSNh8Ugrr65gnun6Pn4
G2ULsejRMRi8RueXGIEQCvZkSlgc4Gp2+AFiMaa0X3yYAtrYaCPhMJjvIyveuvrpQuyYRsgu3K1I
vsSP/ql3DiYwGaWnCth135nFXm7t1Yz7uRUKg+gwE9nJkDIcQ3iLmkSgH4Q9qevrRMsfdVc6XOJd
UgUloCxjfupvRImO8o5cQ9u+q5i5FxFxY+rkWGF/h2g93ttYto3kxnvumGb07jAAah5DhMsMhLPS
z6/SizK9EhgVrHOzlgXCqBKFG1TZpahlK+fMrSRPqTQEJGHJ8NaVqNs8d1yQq1+MOPV+5/SImYHv
sIJw1mmfSXTZSsUnHlciEuY3q+UH7pjyfWtBiKgRhFQfwYLqLHIK3OvtmVV8/z1M5TwwP9uJhPIK
NjMrAZGbD2yIMMPzy/oUC7GE23QGMlp0H5f701tTuxvJUt2ILGi7CHEXXWHIvt+Btm0xTnVhhrs/
XlCdOWdF4mtrVGq0C8eojmF55A1tAzKghbuTvN4FZNTNnGVpGE3J0Aa7vvc+vXLOayHGUBHFEnlp
ZLNUixbmAghrKdZLb1ddScRh4QoquIPOVU+PzZ1rOfeo/+rSMSK2VbmoK2rtyryKe19gV5OZFfeF
fbri83khKz97swSgxi455p8QeAekLyF6kWsNhF7PS8GlpaXPpt5CqZSdZbvgS32E1h02JALS2ZkE
j2W1wfNXx3XNt9DYMI3onNsCFHBNgPz9dBJobhmP/FkgR8QeDfc3AD7++LoxbzC0vFu3nemAaP7I
/ayT1rQA+TrIhjEnzV0EVJL7qzhUU9L+rjVBY6c+yhbuFsTFfouC05G+hyeQRn5Fh8IObJ1qbKkZ
k6WQ95FfM+29x1ZgZxIeMmyLcXC2ZA7F3Cwi+By8QrR1iXG75URyZSROuL9KtfJj7Imx0KROeXzX
6k0cVop1CHeCShkFWiaRzOJD1KJnqEgbYgNfPmmqSdzh61Wv/UA4rJSdtCljC7JaSD17wkwQ52fR
otGaeZMEr+LUYxuqVgjbVPCfq+8Zxy9c8dbBGM+D7ANEm+8rnc0/9QkR2VrAqiUuXt+AXgmWWEde
Y6mifEyo8PfOypgcI4Sr7h6Gk5ZBA9wZoeRzFv5l0B85tdoJM0zRv61EEczXf5MXvoTvCMnk5CMf
RLRzpwBIoFUCWUti0tdS0LUCg9r0aV/4H6XprgcJSuA+k8AHcAthYd0qBQRh4eNw66RsdXAJdBxx
yMrnS/feM+HnPX71IbHGZjcO2+BSvNruYqqqforN1MgJ7OOLwIbs7rTY7DIRx0UO194RO9WtGgnn
nV3VZOMZ0WAlzcgJTW4/GwMvrZ827g4W52RdEZIhWLiVhfhaC0tN5iogmCh6Ey1e4ND6rSQoAsdk
qM7sXZ7Q1QqCZqZytYcNJR0xogjsZ50WMH/j1eAzACvNAq9ThX6rrO/pgTnqIZAmpYONeBsf8ZfG
Ij2hCWTA6uwLodplRNjbjpuEiFZ8XFCOgJ/cXi1eN96yzQ5vn3t0t7McaPYqugt9t7ODeaFcuJqx
bv6lkOpPjf2eg3pdd+5Os1zWc6kaOAgEAiKkYEirr9qGAfFiQVpkEzkMxTbQohU2L6E7yDmzvhLW
svRash5wkvan0No/DxGzEsusEQRdpv8Ee+sTpsz6LT9cA0+BX3xqhkFV/8e8BdMrkpEEkSiGc3VC
RtsX5WPCaDUxym+bhsIK7+55QC487xgtnVWFLRsCAOlPpGaugcsgTVRCB5Exmpd0DjLVpHY2c/Il
RDhdsN+MeBXQcKoktB0BQUhVf600F40PpLl/ng3TykTPSJ655fyz5yH76Bj8NGFSTzS0qg8WSM2v
dGRRE+Qg+dlfP5c5A1a9KTlu8GhHL1NlAXdlG4qqFo0MnyatsNiHrHkJEFcllvxsBuWRQ7jMaAz4
l6mw3qcxrrMQxUjVzg+0CY2nJFQkR4edrSVMHCwCBMkeQKZSBpZED0l6K9D4JKL2ccSlen3RSMPQ
5cp6OLpLkvpEi2GE/zzzJ92nEGZ24H24xfI3LU/JoIXiTL28d37lFHN2LDvitHW+mA3Dp3xsSHgC
wTopGwVQCHJU74z2t2oDD835xgJU0xXt+aSeY4its+vBW+kFVTlgdlpzNa6qswq6IAa92Ih5YJZt
iioCdURfe1rnKcrpQS2g3Ftl3bAmnqCwq77BFt5XKlxa0h/nWBG/XFile288hMCtes94oG3HdlmV
yTlwHtKvfgp6UVqw/IOaOUsMQ0Q+TjwLQZARtXQNSllGZcceVRMfh9XGLoYvM1GNk/szSMS2S6rK
D2NjE+OloEHSJLGNqz21sri2oqhQGPV8YlLSsNuSvJoy4+5lsIHgEHeEbSntc98iMjgNvlF4h5A6
0ufcSDUgH0Wr8RGS5gjk17VCET6y/Waj8Xu7CX9mZ0VpELo4BSNDSq2uLnaqPAA3XP47vxU/A2fn
SMTFC0XzU4Fk7Eqk6nQkf4+QVEaJzSa4asnwQI3RiPLeRwNCgZY8SELLVXM+077fY/izJhEVf/Gh
TLGQh5uZ+oJHmsS3+G47uqgRWpvBG0DMV4GaKVRpEJpj+zv0LvEgEHwoy5BPjxASNzYcBCfGFE0J
21DRH0r4CRjA9QQ5iQ+KOmUiGKjPVulmzW3lRo29BoOxSnKk9UsjmlO+cW9PP8AxTU9/SFITYp4m
oWVGBPFkyRdtH4qHmsz5BNsxOjzYJWBiWDdXGGkdJDGG2WHOo/tHm/GCUTjD+epV3PogFGHUSo0z
FX+PmCF7vas7h1y8uYLihwXPNvgY7RYdxV7N6uS1asvLlI+sd4XqbIGiyJg696Y7gxDOn8MUyRnw
vwQUal8drxmvqZ+nQClZiwV+YcKigzeTsAYsH/BEREfUYfH1yAALh92oxqPsyn0fJKdtW+M+IZfB
KmQ3ds2J06OdZxKhKnrYZKeZKrW3gCodz3SjylZ9ruFHHN1ia3KMG/K6m1TnxQixQ5ykRPC9XPRR
SE6Jbop9t9ZiV+Q2mFZMMyUKbG4eLZVaQ4UWstZhuDw+t5lh7FZy9sHnzu9LpGtDVwQ2KGDII8e5
FSKilhAfTWazvYIQlZw+sox0BaUyn0Wmv7y4Ycc5m+GLVihIQVe+wt+cV/ldXVozQYHQbpx7ZSqa
NIb+l2Vj4ojf9mKNoCWk6JkIY5VDU3J+LdPElnhvxfjRL9JGUR+EuHzrbi00/jVpVtkYRQFT+MNh
BjUfY0insyqOqDGuNvLFKrDoLVsLYNJfxOgr3aZ5IG7QPnFXzdbmLNSnekI4o1nn5Q/9rQJStNDw
z66e87nrOvC1mgSNv+9r8YOSi6OFeHeH3pcl5DmiA7kDJ6hBYd9BckqHsNJf62Zj9t8+mwxX2Oy1
QJdhESlH6qBgPHGh5Ntom2j3s9ye4t8QEhWSmmlMWeXqO+Misv7ZIr/9kPNUIZHMb5Of98u5/79j
BaOw/WzlFGvEQyF4cCiP2VA+QJbLTMouxdWNMSihHDaCGeJp3eTQDW72CbDj9oAfYhzrMvzoE2xN
qznDlxR2VHALLo677R5XjFm8vPgiuHDk4SrstQgFeMRvGGFETUlyyXSHSQB388kBobBsrIybz2Q2
xWop2WjF5L8+Uy4hfAY0X0NNZRnfiRebGzZSo0AuokmAGtxLa2UaQbhVD+dcXS1QaV8zHdze+9qa
g/02jpQghVobmSx7AzZcPHC1GZI68n9RvgJli61xbmJPshd2UUNdM0BwaFRi1r7z0IZDRHUgCCko
PkiTAPWujb4K9mtUCyLw+aWusLCZdj+tL9kSwmcgcY0LtXgeSSywA4piwjmTnBLJSXaV29D0+3Qz
3egucT6IDqL3puyf5K6zPTxO77N4fdGxev932tjyiHVHkGtmcnwUL6TK8mqtF/iXmD1fJ+hehyVd
bT4clA9sj9Ng7CNyHswoU3ynEH1Bn31nLol0289jytSRHLbHbJyn1U6ixgdETCRZEr26HVrN5tWS
c8DesPNU8/SFVXV2D8zhSKbrXeXd8Sw4dL/N4EtEpL8P7UXQhzTgq8BKrsqZkFxszTqQaDNSab/X
3mqQvGSp3xZ2WZQxKLOAJ+EO1cPmj0Gp5TgmLuPClSj3W3/3/2sWT4njaGra+k/aYecU1mkfNpJy
RGwGkgEQhMOXKYN/MKc8cVI2G2tgWrIo3uPVLSCqBHTTT7bZevKgYkcGnAJGr6gxDf2dBhmp/ebZ
0UBE8w3iDbdUawqfJAbgtL9BTSOCLmIw0Xxi8vcjTECwC5WqkmgNf29VnASShzFzlhT+2vbbiF/a
jCNMhM3KWM+GLg1Qzf6PMdGwb8lNYkRuAehZwyEyNew11cVwgLLMOKotz8jRhhuKMf52z22szlYW
KHFmtJ4sAYzEbg6DJZ+TFYpPeth68HYM/dXcp3PC8TzknYsU+AWFjyhR+ilQcs0tx3J1j4FoLvsI
1qdH5Vp5kFUS6B49NWH/PZLcBIjRqL2AJuGZuls31riR8mIkokVPmWQGcBn3gpWy45soLgrlxVPZ
l4mRpF6Ej9vfQmCShKIcSRN6D1dGlwucAo0KkLz1EvoJOflBW8wXYUb3DxAMw1EvNUTdma6/Af+w
fR2lAqRJCpXlg095EZ3dMC6uXG/co5p4j3m28/cC3xiM/VVz65RibUxOOGzpn+9RxQpZD/UqaTbN
NNvrdHKzCZO1KxzZ6u1zo0h3iXbG9Ky3wstumCfuyW2fDTDMv13LoTZxJcEYilyScjZ77htMMM0i
38Qv51Tetb97IMr1mivh872B9Hsip6dd6AffF0o6gliVCzcMrkXDA6SOEQCpry6edBzUBBQnz6dx
Dgss8ZsYaErRh+ZukLSJXs4c47lD+Eo7kUTcibDi43H20LW94RrCqja8EzkpE26Cq7eb8tiS0iVo
uAmr/rlHyzys277xedQcO1AUZ+YhB0L8drW240RMCvGzNAnfGzf3GB7U3N9pUs4b1SvEYES3HZdG
vffVH9f7L0Is293by/akVqYCrUEuBX6sesx7xu9cTadt4TI/5Nw4coob4m4Sl/lByfRy4bnNMwEE
haTykPiOlKnVj0SXmvn2l3yBxtALJclJvRXo0pmpptXS3PLMAP3Cqm+D9s7A/ZxyRJvVnDhIpZIv
xrq2t8yrlKt3/hZ3OM+bbBrBystGzMU6cbycb8WqRhkky03VAHBHS6bCDNFT1ZKhSuF97+CZr6uG
rWsAd1Up5wrO7G69IghBao6JT+p1WmIOzZbXe7e0O+WKc+u4x2UpSdSY6ljaQIn2h3bpCpy1zTEi
BOuN5uDHX/V/JvsfxYKaV0xmYFFcmV2a8JV7yPi9QNf/Pq+2x2DiPAtWA/wDHqL+n3zHTIhzYuFP
Gprln88JeUwVizWZh1jM8fy2F2ZkTp1M6ZijQDU8kV0RsB6TyKr0johRrpzmwjfUjDR0aJaM6kNr
yaHixgc9ae3F+00ac/NWQtUv4eSBJ5eqlTVOyoI0zzuo4GI92yUoqLT5aCFoy5WaDiSjgleZ5jwQ
5MgsZ3CFY54LfU6ev50kZjlGF1CbXPhAhis4tm3NmkZzzkQnZn7980Y+gAb+Qz/wMixzsKmUlDxp
32NeXwFifE7dw53ehaCa0uYihnzPbrgBLKX+ea7CPKa95IhG4qFf71OB8rmGBg3H7Yeb5ylHkLAt
JXOrWHZW2jbR8CIcHYbSkGsvykaQwFOgM0Y/xrY0uwC49rtoSxWLYrD2LZfQ2efbClwz30LOcYQN
M0eQqYgcnMaeqNkLcGPBl6mhnOkU97if4L0C7VGvXGdi9lXfKEbW2+HRlrglPcp5VhK6T5vjVHzs
lyCTEvrlVURExDvnTgCO9UfL2/nB7N+s6tGtfOLyacPledc/wPM0jL8AoEnOqpJBuMaRCeqvLUIO
lmiKyVCnJZJCQOHs9KTg2K3pxo1FF9MNHQf68EH3ZDmHEIzZd+4wdUJxtSmAkxZm2UTuhRnwMhqo
k7Sr43QU5hVzQJipqlugQbnIQcSGEIexzb96j80dk7SBOOvOuTMGtGyQ95nGAkQ9CryTwAMmsm3C
wqvWEu+tnPB7TeMy/2btt7msLtZ66LDYa2qs/fIvoo2XzwLOqTXN1IfYc78s69IvYuS5Zsf13BDC
nFB9UwD+0VkUf/BuRVGQcI6bsee8v63KWn86IpdgK/1bvLFZaHXqap8eJmJXsWzwu5YUft6K6bj8
7AWamXVrFu3b/hWTouokJuhA1TZNssVZR0yq9YOA7XTns0gEGEa+N5dIAmZSNMvP7m1X5KdP3HZA
YdcvXvlL0wiqteR6EV0FmJgpeMma4L9qVLezVU804w3KbGokdhbEgbT8L9kLIcXHWVDENmqBwspX
+U+xHwoZkVRcin3swc8dbTwkNn9APLpLKacL+3SYsZ/GNslt+uyzgFQkysx/8b0+PKo1k8xnb6Jc
CapMQCOIr5of70eK7xrNyziLKeWszSfTeMCB0FZtVOgXqtIyk9S4vqeSvM4b6uM2i6BOWY+V/boV
H/JVmZmtUjG0FFZJRhT4DFHUrTRjmB8Dd8xbFRx2zcF32ccHTo1Le2EroSpIhI+k5loddARXTHPq
LEsXk4iLf2dHYF9DNk+dcZaQ5KljUnqF+E47EUwZER2XS2NWGtArig72+cLzqwufAFbW6rwz20Mx
Gfo8Q3N+XRojXTXmG/6DP+AnPfbwpjZyOXz6WnTkzA0icrK37I2ZtPIiTIat812LoagX+Z1OMiXW
La1oSLVIqj4Ts0xkOaHDCLJAZAB7ZG14zllgibDHoIPBSGzBY30KjAPnFZxAuLg155Z4CEzc+tvd
ovZzprkOwR+HUlY90m4yI7POTW+QAFcuZcXaypW50OdjClPr80s6Pf2kNspGF4us+zDp+Vbb9x9s
dm/n7PVkjB2fMDoken0+NbogKlWxgvp43oZl895nA7CwKfFVVh8CrdznZWusmWhGq+UwJZx0iGbL
xtJA8N25ecu6/1XegRYh34Ovl5zo/7/sc5xCVV8dZml5JQJMkxt1RRjose7lEM85lL5X5r1Vue4Y
CtqpDI2LJehbVZHmdH+ecWtBLeFPm4qzr64RAntylNM+dByZo79tkLub7glvPC60aRVgZb15k9Gb
67yaXWWgBlb3689c5zcj4BSGY1XsxTiUT7aPUZJqXTlzk6JZbiYpCl13I/9PftrCn1SuIUMd3G55
zOzb5gCMpBC1HRep41ZCHittFWIeL+U1TgDu7TbSY6krfskYFKriuz3cfycC+/Y68mldazDl6jxy
9ynul6Ha0RVRYk/Xjn0E2xEzw9f3Z2vezr97DAlTW7X4kFan18Er9VAM3XhhROG2KwZH0vep+nGy
SJYm0znGukG0GHiArg6lwuHDljBve7uVqDKUbTzlB4bGQJ51VABDW4pXzbJJiv69mavAyOGprvHs
FZCIw2ALxhA9hRBAzlSIXeaDuOndLeZP5x2nwiORdw0HIy+6pk9s7etKWnCYAqwyKH/3NTtalU2+
9JQhkIMf56UVYrDCaPA4b5iwz/O9IDI/CpSlIYAkSvDfF+LeeQNuOg+EDV32OWBlgBXV0LxzFLJU
pQZNUlSsmwuDSE4+Kx0xuAqvcnbEEGa9jzwUDJw+mJXY7NxnrQW/qEbzZ3S94mei4nkRNGF86Xi5
qcCrWasTQo+uecU1vYVHBtLOds8fe/BymRuA6Kwj8Zscx04I6E4OnGmWBOCAwezRcsDYtNgr23ne
driaFcmygY/O8lVBpK491DWfkjvWY4oU3YqqZDt+Dk3ScWN0rT2TbIb9oZTEnNo1+IAFAPMEqE7H
RWZwLZAs1rcTzsM9PcZAvPg04oG3JMk2ou0jKXakxv+Ap2+CxZPumZElxz+88Beas3JLe0XWrdwp
EG2s3mtpjcIey9AxI4b7LCjCOU+6eLgyzB8oDRL1kjU19jVI3FsoZ75qH1DCPR+Dz+z8QARNyUxj
IG/445Oedyg9xn91FewpkCZlceBczdrFu3jWYu5A3Wohd3XLKgdogf5reYS+XahIbUK2UIQz2Rw8
WitUp19wMspIuQLiTKRfwhX5Ii8l+KTqveTBNtWyO/53WdHntWNwnGYXhHfjNjLehl0VQF8jdggW
mmn9ds5K4YcEhmfoYMMOpLDu/uHU8rMJy23elPJAlk6iQRpUd/R91Rn1emHWg98k7wQA4oIW64nF
cMCAGd8MehATxtUPcTLihFCmQiqO+Nw4eHPO4QxsXFrMka3jkOQuyXTizGRfJlNkDYAv4g2/PsHv
C7S8ZIL2kXoZuWolc9KU+j73FO3uTYDP74WsRf+vdlmwCfx3rWjnDCJXqLXd75Tp439MLY2yikbD
izJCgLJfpeMRJBEsiMgnjPp6l/7mbLT3nidK0l2lWIKVfOyHEudIjIERuG6i6oyuhvVC1Al3cDIo
u6OZQoomKnAEuRLHmQS3cxQzJhh2bkrU/d+cesO43o9iuZg7tkaVBxDx6KPkKLxbpChFENsOq4WB
yRd/RQo6HT4ZzbPVr890V4U0VL2o9/eoD4AxDpcrVCYQLceEbpo1QDhiMed5+cQzlHBO06Nhh8Yn
mTvDnTpvplmF+HrgQKcjGIyG6US5XUVFOKg3RdrYzsWhC0XwVgW1pXQGP9n9ESWnmtLlM+zMZSR5
VM7XF4AK9M14Z9beJDfbytm3nLhITN/bz3WvZ32JeyhxQ+AQR2UNX+jQhV8ik8IzrVyhYUTbGN32
d69wCLuHpiBzK4KYbLBHYIpIggSwMo+w8AQpz+zPkqK0Ye51VIt1nd4Juriwqym9Dee8fBdOPLHY
bUZH7N+jvZRNJb0MgcHcMAT5CZACkss0KpTuAiTgCERTgYEu2XcGfmlPoLHDtznI8ZisDQ9GIL2/
25c6lvH4TFogi2Yhg76gzriZG515KtxK98BuErGL6+My7YC7rXZwM6dcOPafG0Ij++tn6ecF1ZUB
qXjx3gomJnKuk+L/QAtjcd3YHdN6amuw1X34KFRs5s/6wkygmZsJxGXQewGh3jxyBISy+kk4ytae
6sMxn2Vhw5Vx+/QfTu1GyIG/7MS2uS1EsyMgFGQ1TsKtRwYsaWc39xDVfx8KOynjAy1WHo0SqAM5
aGaad0EeekRS17JIXIgidh51nkELjFk8DePIvNcpoc7TMBV34QWvaFNZkVw2Jxbx5V/YD50Z4Woq
Fi9hzefq9bNPQJ2dBFK1ZFtXOmqGy4/bIJgCI8BKSAF4kZZZB3jLFiWhjm76YEFu7mFTSi7+5QB7
ZN9PLtQmTu7pLiULR4PE571v9dju6bwTcOr2JnucB0ha9oVYQLk6baraytCekdQap/A3CwVS8Pgu
icZkUJk2iW3re2foS4DouP4OxlYvxfR7FkxVLTyfOQr8T2/FKE2qAo8AQlIKj1+Ci/pQwvzhLvM0
alZotJ2ue0qH1p1i093wkW1ccDY2+wieEgCo213MziJ+xMnSKnxuVqGqlry/PUu/VrVqMJ6Iy+S+
U9srJ6k032A4BJrp0Z1x4adX3xA/A2BBrcTiYLZXqtBj1qbvzZx2WAryjh+4JMWe45FF7shVR3bE
SUsSyMlnk+Nm9RdBA0Fqb4R2YW9AR6DP2EoNfjBSx8nK1ywYLX7izWU6KMp+rKAWRPND6mYdVcH5
i9GlPpKJzk2AkFCpZr+pezHah+weknHZSJ0yZkl0eqw2q5YlVmV+drZZpdo15d6wCw9HZ5SnC3US
Ymz6VBtKEDzyrJh6UcyStP5CVijbmtO/cZMy1RcPht7+c/5+HdVkyknknlOBzA8RlrLm43ikPGCV
8dfpZLrzWGC/GwWgas5wpduYh3ypHnQcjA2KvdamNVc3tcokuh0eMm/Joa118v9wzz3XwMTnd4j0
451sgFsytRp6VCQO2peXn3Zh+RHKrS5+xg43JOCvFYqV9FMsnYY4AWXTkuml6xUECo6L/xz+kNsv
rR9ZL+qVzVuACNV3EuBCpxUgPXNIemBNII7lVHzm+cP3B03fuDXY+U5W3YGedX2ogXfpymsMCcEu
BGvJ7XlJWRFLO7gRFwHEbQukXu1ts/oeN4d+og/hJywXcMgoVc7ervR0ucN7Qyow/tSlEFcmaP4l
oPqzomyvjvSE74qTWvEu2Vqo0L9oA2GBeqIKrDpMUKH39tltbybfIF5dwM63RWZtstI0xKck75dW
on4xHZGQrnkCDfhQ8zBBwgybhiRoEVkmDnaZex0F4j92Ect1fp8vvLJ647qJYhxwVh+u4ZzzpHbg
q427gTpMqIMRcbuxh3I3nGczaD6HFnGELfQwhiIB+Z129EkhKZWHV0QwgQYgBZJbcRPVtyA/RQVg
jrAvAE1rIM0On9lvIqnGPFODpDFa1nfu+ehMSR/Ws6n1X0QY4nVUf0NSIgFkToOn8ACKr8pNG7Rk
G1wTiu7utzJq9iRaat7X4HEGAA4Rz4RZi3vlpLWh/E2j3GDENg45VAZkubboeRuNUKSfT5Ri/I4i
uhtBpZCWP9W0LkXQN/HUAvgYQr3KTa/mtqmrc/5HqksWm6zQbNj8n2JIXQil8AzNfGrwO/5PNlOJ
Me1TK8mVGwMAy0P2GLKCUiUJgzgwsh6X7ykhmEpfFpKqZzk+PO8NpOy/CjQP2WhAiiDfJ6U04RM8
9V7muHMydyBTeixyVGbMgQ63Izp+/6KUSiaZTl8Rs+7M3vRjOYeuWf2apUM6XKbo7jKPszYGyiZx
LX8VIA1qvft2Z6AocG3nm42Sjn0DAmKtxl/ehcZRrziL02cYVVNXPvV6CdsUOuUb9PF65iolL8Cw
cOwwfZuDY9JPKLwxiwI8/bgACfaTVgP7lGUAIl+fZi7Wh8vcZJH3dYvgsWxRlI5iqB4CNj3oMMO8
aAGDvVW/9JfDUMqsVQQtE1amUEtOBWcUBpXkghuYPj3ovQ/lZmG9SgpXBCNg7hsROzBkZ0TgU5CF
6UrhisByf1Q5O5NNvC+OLSpM7diwnl5n1IAf/eS1o402oKffoxgAMND0Q6JLxqZ/aLDGg6sXS33Z
bVU7YrlbjjVyUSbpB/L0ZxFTdkOSsFAxWBQ65r1qMq67Gq3Hjtul2DTacjDbvBe2ReGq4iRxVILL
Ctia8N6eSB4AAbLS7c0OIL+sJNmkNCpvlIIpYvumgTvQ4De4WMBfnqY7yBZOh4nldyAQXU01XAdw
hELXv0vdtl6rx+b57fYwGxaIWJKBKCHXL1fPof+XzS4uUxhVIPpys+W1DS5uZV4shijtlQRP72ZV
JbZj/gbLYXOoyiY55074V1V1SjMrpsNA+Wwn2T2wMGOHmmay281MSE4M7b+9u+kMp9SGzuY6/6Zt
dfR+LejpHicVHIg/upkeYU8jEN8q5SVyPYl3LZM/G9Bo9VDPIWsLgagQ5oobhAN/I7/Ju3q/YTc1
9ZoNcYcRbT5tv/uwETUTfvUrZRbGVwdNlYoCLjv2/8ryj3Rcrut/yjN0brbIk/6MUdguSpeQ0Uel
3mjGpTyeI3aIQ1r6XvTiK/WJVHcBCDnu2vrcaJ4hOOokyCVZ1wEhqfax3w9gljXC6ZZ8Rj3t+A/i
nurccVz8xZWdbIljwunom/636uVT+sMVTg2ZbKInWH9qHHUg96n72AU4iYoy2Skb+Kr7Cm1nkBKJ
4kY/mQJuBWBWZY8Rt5J8X+WOwderA//afAP0mbJS1yqjFTHMCUyUqs2/NjywKVbFoiZGj+cbaPQj
RXglZqmYt7FQzO6nnoD51GCxEGUTieWb8B0UMqAq1zrFpvMj9cYQDcj5Uk+4jderx0WewAE9jU8T
gUn2Icepx9kqmc/qGGdKDBe7NwsugdceQTSFI94cW2YZbzPU8JChjGehyckf08U6D0VM1lR62hEc
KT8QPL9FRjN4oFbPM5m+FwR/zfMw0if76V0AGWfgOXYRm2P5gNV7SM94u9jYzSyBKgmXC1uQlrDy
josFO+5SY5KlBviKf01dd/WMJWUbYiwHoDCYyM6+kQ74GKL1t9MI3VY7AOjJFOMxt76Lfz0FLDr0
HS+hw5zfxtNlycAg4mK9dBEujTjRu18anoxRiey+hrQVDWeAwXzm/bwsAuYZGZ2paeojj1wynXJs
5d40YNVLGJ6F3/ACkn+hix/tTjWxIZ6NxN9C5NWIWGdG9vreLCukTolwLrd6vtedaT+8XtYVKeOs
4nfSi9om/pB/mD/eq+6LPBAgIRKu+xkZJkDZicGac0BWZ9+JDz3k4o6TcziO1CI/uAD9jcfGktp7
x+oWLozhPnAkLp2fy0oBIPB9I2zZ456HyYSAvOCjf88MBei13vqQD8NFIYD35owD7gazWPdUl/2h
KK/Y1QwchWPCA98xDYHXJaSEitxAlpM/ecCM0LSuGBjdTGxASWXpw6ncOmtRRgtGAoUQ33huSHJA
8kI3zWX5umIDmYVVq3Se1C9I70bozUuPWEIxSiyYcHfgz7tY97d13wiwUbs6Odf5jL6/Nt3q4evu
0A50+lZQQUICl7d8TOE5YcU5u9fhXUZRgx34y7REA7m77o5fJR24juAF2Zmyhfe52iPU50j+qDyr
9M9LPhvsbu8mPnimFYbujFFojbcMW82Yezw8YNnmEfAhiuqIgCwG1IBr3rwV5U+iFZF7eiP9L9Q0
gjSHWiq6vx3pSQmCy1UQ/i43gWArKz/eHc15PGRG/wMXTWA+UA31WgrK3RPHQxsyQGdnyfqwI8pP
wuTyH6Vxd/3+M2TBkrmCQm9KsomvBRF9v7iXOT7sYCU/E7kZbu6LnsJQDdqU36qWfAU655RNc2JI
HWJY9Z1vqd3xKadQW8wF5IOyj6hPv7pBRZM5MzRGyWzs19o8+/vAgaBH9cMUIaa9YiLqbcVqzHgr
A2JlaAbBUzx8FglqYCCAsPJExZLUs8XSZzKxidrzR9pmcBI5Y9JrzVS4FCp+BGbNE3EsL3Blv4AE
f+GBdeWVd+pLnkQjA16Pc27FmXqiZBIbcqI3GMDjjrXH6FnTLMWI34uB331GbgE40Hvxw/RFE1Tr
lrLSnwc4CL25PVFBlWNG4sTJU1x6NZYX7Y9nW36wsttfRcNn1yZ9oVK6G1qamVhBu6GciOi7404L
3589EWjXjFPIRhHExoS4hdiFgqTqmkfxn0gaMp4B6VmMV6PifrAJWzo81rdUToWhyu5mkOARzVx9
DmDtWJi4DZXYvqxx+/xd7ME8LRSjH8tuO8s2p+/4MK4MgU0fBoE+7KeneKv+fSZ5Mlx7wety/zDw
9FHWoIuWUhhICM1J9viV49TyCHh568G5a9OTA98nTsArYlJYDnQZ2n2b7I5OPCxgmBmfNA/iUTuT
MckPWtpSh3r6gQDJLMT56Q0OLM59MO3tGsyqkugtXWSj+oDBzajcWHVlOn37UVoX36304Lh50JeA
bKD/WQPEri6OrvLg1AlP6YJACvBN0nhjehTuMSu8ZwCv1zQR+EBGHSLIw2j0ZsOjX5TK/phkkliT
48nXuj6ZTSWd8Z2xG8i1l1QjKU54gLPVNE0sHAccWPcsxyqKt8zH7PXpylrHbsMBVi4z7qOS2tLn
hB02LQENnMyXv3v9NiAPfxe3QoC8Aj4chWlf2g068cgq7bRBuijLJUaPAa6Th0SNf9aE4GbmE3fR
W8tsRFlbECryLQkPBAH6MOh+V5k4VPvWXz1IcgzhuYsdl9BwL1J2C4hUbkVLsWhq7/1K1fhQgBIz
T07Etr1+y/iRObiCUsRG9mTv5j5mlXCbg3mCXK5/3+cVEVnkgiLjI+qXDP2lSI6GCgjW9lyY79SW
THMmRaIjsqlJTGV25oBpmpoJ5ZK5aoDVtOKLhOkm8p+FKb1u+b8IwlSACbPlwLtH7BsTdlARZEMw
9cEn39vlWyGgGC7wK7flEURF+QEzYLlRk755FsolYtNqgfY4ulIJwLR2md6j/K51oktJYNLNSQKk
ZvOSvyFE2AwvHLzmAdh/6/HncAfjq2H5vtfvzKShbicet9HaC7gC/tlT+UFHrZYzcMNN+INTyV2Z
60WYYAWoaGOWv2wT3XEKMUgY4Xuq/SW4VrMZ2fGWaSGv/CxcxTEvRBWf48nmmNVobwyIp33Os7b3
kHTJNTU/+5uMEMKVuv2KGyt4LSyFN3xE/cRd2fGZR9/Wiiw4rq/rUNwul25LVqUwjj1zXBL7HmzU
2CxD9fxJ0c1XK6fq7BbmJ/zu9K6bH3op3wxGHlEA1tXurr72nGIcFb08gLXkR283KBn82hjScXPe
UeSn1a3VoHknXM77eeK5Jc2CRTNNT6bky2PhGKVWGujWH/7SSqRyifui2qDKajjSnCsNZbkCbApY
X91Z29l19lHVnXgP2g1YPEwZcsD5IuhWfjM+dyo0QsgdvFR/aBjGzlyZWiavTtfclqotiTCx4ovS
BoEry9eFoZS4R4oObuY518lK0PXGJWlG+7j1Tww+S/rARDRzuDwAcnUsb2z6CZdMPdKKIjLTIH5M
e4CuR106kZKhhy0SjB7Lo8/7K2bZV43Kz7zxiqYvd0fDytilQ3oj8RoOKKiLTACBcO3+feG34KX0
slRRKh+xOK2Z4ABmzY9O76FvSxw240Csca8tYvpfzgqMsTRjYngqtZ3Nu8C3GAsSSAwAHDaMqbkp
uQVC4kgVSv9NTOPiVQrT8JMdWALa9u0TfbTzSHkRXs7lAyy0AmUCGJLIluxblTLCao306x1GinSi
ddMZIbcSAVl1o6BbUV0rgM2VBFfBiqWC/QVgLwBiq/Z0iFjis7WFQkOBhEf4jYXOXHo0Fpdft5lh
Rc6jTo4MPiUFK3z3aPY3ceRDXKXfd3vzW7soPDbti3E6XEqQ+a//C5SygEDbYpfTmVl96nw8ZC3y
+Tb7yi8CK/lQQ1kRWvzwAGR0HczX0qSIL/a2SSeXpvlCrlnUhmUwhOgHgeR6W03JvgPCcY59jzIa
DeF8ONTGNWn0otbdiQM5TcIH/R/BBT5thpOXVumOD6gyh2GNPaO8hYmmcG0zd69dYPWy72NOjv33
IeuJN/8zkRWoznmmtnCXg7CtRcGuOGVBD5NvoIRpH2ygH5YJ+kfkty2amiSLXDWnYNd/gh7LsCFG
pZvPi8dyW38BxuQmxfacSvOI1vKr1rlhYa14pPXvHoRDwF4NZLV3/V/Wuzuf+3FXs5FU9+nNjhzU
J3kL/0AzJIaq3lHq2hH3KOcylpc/Lv4YOphsr0WezXALp4OpT/dKIYzo88XBTq/hqj8UaiEeAPhm
C6Vsk3P/FB0FUTpYFTEn63fMZ6W0bpRB31czlohJtNZFH1/Mtsy/X1vUfp85G89BJfAYTmk6bMjt
aCYHK0C4RW0m+WnXGjT1QoukOyYyZgZy2sqfx0ZO6pZ0as/roVjGxW+GTDSCm/q3Bdx1AYyqoJK5
badElO4NSglofE/sd8POnmq+jvh2NYRzOTvJtruMsYUGQJJqCQn/VTl+pfdD2ReyS6pSZhyohpET
rKx92+ROV5bxkMhg7v1pCtMq3irNr1ZvqUtCWdehD+RDdLmcHU43I+DFiWLIfqUlmDoCoACZkm81
bu7yQVJNMIIIOm2kDJeKQClR2REKrHQgk9bIVVl4wHdxxvhYNiUpnZpdBXJRmJGENx9PsT69vUjS
MDacr9svrFqRN0AQWjTkv8MtWk7r0CeQeYNzD4se02Qg3TMlXLr9JsemgLb2RySVrOalyIMAcfaH
GIhD/qHmQvK8WHHajJM7G/j8P4G9vcqHuk8T/fbqTeQKc2VFVoAhVDN3Am2peCIesItZjUnoWaJZ
ziTyhEyxjkrbnY7yzLq4bQOW7GA6FOUuFeAQZI5seQ4TMSU71E8EV4hORIgK/MtyF70G+Rr0fj/p
2oX4SAKJ6t04+FrICrMhtr/cczs2MrC6tmmfJiBg0tlPoCGmcFBeDHud3VyrzSmtybl4N9SieXY+
hpfWgYLeVRw0omzhEadfsSvfsEARBqlrJe/y8jCsA2bWvLF0pwfUmAoE2U/xkPrdjGFcfRuchiAq
6QX/q3vMctynjbI1REJaX3Y3NbetwW18fJ/lhXTgjFTViwKAuKSLIz46Tl2W5xrufKwqkgh6hWG4
n9HKwl6uD+ZZ0ghwXfCWLFgv+4cnbh8eb3B9NdecoCMUq9qSQQgTvoOlucmd3SEBl22rp9w8hGtO
KvSf+FoPC35eAhJzn60uhTKMKKs6dnRQmTwUuhP1+xQUxeDSadYFfpDJLyTFTCANdsyYZTnAmffK
saOL16pUUsoGJwogCczxSy6cLZsNzFrctIMqmmSdHS/m9SIME6KLCGF9qKlk5o3qoroBryVcHOGi
u/0/yZ7BqNEsOkP6atCy3h/xix24PwT3/Fo90hi+EMkWhspmBrGtiSsBRk7NRqqpDZfMl4+ACf8M
TftxKeoz2jG4rH44UK/N/6WpAWF19yiNThUcYjV1Np0/2JWdEokmM5/HxlG9gKV/sIz4EmSnyzYA
eLAy0ixf90Sc1fr6EAliax9C1vDn10IBH4WQggnDHJTRbdo13HIyY93fG0naMtjw4GTvLzZvxwPG
0l/gfi7HjQIsfqfTljGkU9ZzpAY5tRCv3T5hVpezTw/FgnGOQQF5M9CJgW1ZQMz+Qq1CkylIlTnX
pyYFYS/lnTo/25qf2cr9c5jnzj9OnpAqttHiqikvtfgHl0XCAUkl3X2zFnh1g9NwRIMgD9AXjYe4
DXfc4irao/CasMUJxtlkae0DljlT6Z1Wo9ZJAqa2tZJwPTTjUZOZwxxkutzt9yk8LAM9OeqzyqcH
1Oo8P6U7G7imnRBFnLmB6k3XaImjnShu+owyY6V/EmF2zS4Gp2V1WcgaExrnI90seHrocgvfDmtq
BYw/WGdCWX056LDVT/qYd/XsxInTMAZvU6pYQw1PqJmjxcAXKYK5/0O1LJnIIFzszdcPhD0D850B
L7y5FXz7ny0HryFDYzYWKtANSSbRb84N64WFqhNIa3k3DuAOfPiYMxOXJYoV0wU67sKi1s0hAphE
eOQrDjGCD6dLgrV9WdxbTlhr5QGE0iTuvxsWHqswLLEN9fmBJ0tUT/JfyufvSwxgYFfuzxH6UEJJ
et5ee9RopY7LXsT05FceTUdR9bH6zd/XVqhfqUMxgDP7lTgIHHpAydeko2IUl4PCj6wBpJV41fnY
em6658UqUadvY74k2ApuW3UbC0ssjlll+jMHH73hGr7X3qdqDW7x7iuG+YCyoDlk0pmJkTQkL6F0
gzkacbTyH5Q1Ouk0flH4bbAFGhIlMQvS7RcbCW/7kauC4X/0frFnn8DVi8tZw0oc9pGiqFXB8TMI
qFiPcoet/MumdkXbTbTrYMoR+DUC1+UKm75q1FcCUVt8+UhakG21SiwS7Lb4H2i3Bt61u/UnbFI4
Zu1jj1RoFfrdBZVWATu0L8wxG7mxsgqRGytnk4BkaL7lUsM8AwQLhVfwhDV7TJDYC+DfcyqJGxRc
0Uvf9GP1EpoQZxmLFvhyyXWxHbs80cdBykj7eMfwuuM2EyUs8Kis5JChRDStKuOeO+awx/FVWtQl
vM5SZxF1sf0LZeF0Dkqf/bxfhGv+32RYxyUsgbBlMRAnAH7wkOqjCJFo/5RQweIScRpJSCN1rMJF
Pa0cWO0O3jpzmPSY6M+SpkB3XHwzHGH4YtaVMO+h7Sjz3ehiAVEf5mUWFKOzLuUrorFxurQzbIS1
XvrWHQvsFNS4xP2zMO/odwEXPeJ/Jwxmb8QVeyTfMr9DXj9MGGqmB89r+JxLt63ACFSIv/LMwUK8
6vvMXR0gur4V9KgONfk7QF1xu2KcJwoXRt/aWf6szbTOSncWx4/AGaavubMV3500mqxdzzzpaGqz
jQJmb43WJ1AT0/xnHFIhOr8WVDrDfmA9Nw7TIuFXvQPZGgSPpxMtxWraC/vqr+r3ntAFZPYjIvSE
KGQ1AVkYrH0GCnO4PRRjGTs+roAyDXKbjqQx9RWdTGpFhgpQKKQSPz83jyfG7A3MamVdRSyrsmPy
/cf7B7EDBv+8nxEYVzLLf19cPs1k6M+jOv2nepvg+U5b8QlSDwApW/hZ80VxZSP9Xk5OXrq5eLff
UXL7WFkrARH+PefGKQYXS4pHeonuMrypa2w78GoLCCMlmsqC0U4jaKb5tCkc1+kr1Zu0C6XmxEJB
SMZDeTb0fUAIYBlIiCbFYpGrMXsrzWx29VEj8usBCqnRGZmQ737YJxGZqk/MZKDmh9FIgDMDU020
BhX+qa3QcC0w1xqUknuEjgtjp8PiQz1qBMFpYuVlm4jPhFQ9cQDvTzWTJgx3cu1eI5HB9HA4aPK5
5E3It2HDW/pp66NPhRnPU8rqYdiiaMUexUe0aRRIYQYdBQv3PJ4A325qMwoltZqNWEYt9jwer6n/
Fqy3oq7NKzORATJdk/Nb6XKbdSeF9QA3j215BIUsDPgvrJURdKJI506hUJRxytSNoU3vPWS2hz/u
lI2DzzbA0rhn8dEhpW3+QvamcRY/uL5MxA/0qYjqNl1RK+tyss8ZT41KSpXMLzn+7es+Usk3HkHU
9P9ru5RFxxyGiUGMJg7U5wQcLwwjDfqnvoBpsd95H+q/aGDyThODpVRenwIVJe9e/IAOOKIk2Xwi
Y859t3mIl5X6MvytZyzwBZQjffTPuddu6YxROd6SmjjjaSmbBrtBSdG/z8MFmtDFmQ9BYGbPKkeC
BH5Zrbb7nYS84eli0LLDFrpdzFBGJc7rU0KIjrvqCAYmUgKwf5vN3hRA4dMQDpXOs0hONDQpRYPE
RZ7WGX2qtIlTy5TpIRn/Q96LkP90ytl4wgEGrnu3uELWfTinYGb4Wd9k750EGV8rV6GGfNYsu1fF
oVtQ0/V1ZrDIa6JygRDXLlBKfZz6gUAjpWUiWa7RmPtsQq06HLf49L4Ml3x2JpqzQjcgzGaSyOHq
ezIk3kauglyLuj60UcM6iSuQ2FfkrohAI3f0tFuwNbR62LM3HGT3BN/a2VnAOuLJw8JYC/4XnPCP
icIq8E1VPTu6OkSIj38eawuOQzDB3++aYxlKW+3Kpdct1DYovflqkeAIryGm5tLMapDW3y30FoEI
wApIqOPw4PEVE8Ul678Qc0//LVeIUmPA6pRM1QmQZRoccxdP1T4i3v3f/XsDEMgn3yz6cqqxztvV
6VekJ5F5gBIoO3/2TVbJaAs7mrkRZx98Hs1CckJD/q/62nY1RnbqItkZWMJiM9GWF9VSU45O/cJ1
d/P+0s5M6ELo5nub9ngJYHLiKDmtsoyVfz49Je2eb9aUVIkB4xBDUG973gYTFW4cSYDP6HwjotUm
AxYemUEx8pmHANYxzXboCi+bayI7r0FZPrJ3ypPhOfIr6l++HASPU6rjSYVhtxcbCdA6IVIyX+Zh
h09w/VubKOO6/xkp01zEgjSxN6HNMczUi+NplNbz9G5mboix2eAQ21kOv1kMpbPIIZMCel/VgF6/
JGNWMpmaPeDZyP1W8UOkoZFFcfq7bIdl0lcCrLwayCzFqKO2itZFj4OzgPhHEAoUE4YlxalwXPR2
NBV/scvq+W5UTxL40fgmznFFFHzAT9LFAVkGWJwTUHp4otbmL29mdun0mP/5zuBRfs0cTmpVQVLg
Cc4NosCrhCcb778I260Gij/zYCRmaQut4Mk4ZX0za6SbRowe2B2GYx5HfR4PUJlkdkd2amUrTecD
z1dOBiTol0nVf1hbDDh0vNMj+VNv7uTy/QsK/yA8KFnvHtG9BlzAeuiA0B+ZOelHs6A9M9cLvD68
UlO+BRrKcVe8ijVw7kC1AnDlAbit9jbcmjLS57HkOXtdLd16WYEVq8/6X4JcwIHt8XM0+Rt7bytf
mo7qxGIGhUPFt0eWlL5QQkoXMtB9ZI4TMVi1PcJNzcGfyi4TrDc26rFsc3cwXIPz8/QQ3XfPT+PV
5vYnL7sBF0RbOvYTEI3lM8LQQk1ckBUyTAqABBEDohqipCItFuXsUgKKAV7/AxfxtKhU1MQo/DYu
DwLn3tkucee5kt3scrWE7KSGPsJyF4PBZjzAP2MukM0WORgIrCjEJrYCFvf3ZSUhTc0IwC84GRF9
9eRqYlnhAM9SG7NI8jWv3RO61IBEfZ+oU/21OqzM2GKles14Q1ZXZfKGndzcU/Jv7ew7oMwnMUCH
SoCKiZZ35DAV2v8Bjv4zExe7NhQafTznT0TIvV/dUB0YcSLn/MU8b/yivezkXIl3mYI/6yv2D8JU
+DtrqHTLsCOd2EjV3ubvb8tOUSJfJx8nonCUuYwjuoxeVf7PdZgNl7+6Yn3qza2JdVY7rKJJe344
Wqu6nOGrXmlL1E6SbebIaEe7np+THm0PJnuvsgyaMVTq1tFgAQn9H8tJyQt1bRz2WlN+S+/UlqyI
tRy4x4RSFsdwIbbgKuOkQu+F39soub0WIoFFENGo14aQF5Nw6Rm+6L3ufj8oI4UkFMZNwd+qpoih
SDCuTi/hL7XMeXIYwpCsOL05qtyI/An+eAF3mJH8gKtURRtRZQOVLrzNLr7tTootkYxa2Py5tmDs
wgw3tZtBdTxuPEzEtY2OBPJZg/R6bxVF96KqODWTAQbTObrhEbBifGO02MMdPzKZtPPPPcDv43e4
aDeBZF2V7qNu4Ct1SLRIM7X8mpG+o+geMAp2FE0VimLWMV5Q973qjUb8v6QminVyLqBEc8k3ykZI
mRfpM8bUizoJ4Mpd82gE9gDT+568tqPo4YaZ/LRDLDDf3RhPm5tzpb/udoIWl1i0Q7T7TPsludlq
iaZ9BoQJy2T8yxLK4xfyzYa5iQpS+90ktLqzo5QsbshwMtvalSORM+TcbrsuP2YlppUs1yZxPrP2
5KaFZ7jJQtNFKBwbAahCXjzfIvJCjqQkZT06mULpPmum9cn4QkVk7apLx0KImDkI2BpdnoTtkA4u
qRH1HLrrBJjw+HyqjSiuQg4MMAfr9qnnWqK5w5UWcXwgr2IAuggy7b/FyuqONRymbLzS3lWIcOlw
FjbTeKldiRVHWwqF//Z8QnBtv0fczD01UyNs5+ij3MeMcCa0mX20iZzz3LyroFcerBWjN5NnlmxH
DdwxyRb88CSN3iJn/ts2E1l4xibW3w/+JLms3K6NdM3ip6w8xWjHPhNGCWSBTNCEuUO3UbS71bpi
uQNDgV50neXG3S5YuQ+k+RRSDA4zqgclE0K3Mn2oNJZV96CftSn2UuBXCw91Dtb2WX3KMpNwyoIn
NXvB5iHWREinl2k17ZDsOdigmu8pJsVsh7ofFh2OAFnKjYUcuFrk23iQMmIrtD2HEGnRFBiDnxO3
ljVQUqZWQfnC8b2ZkN2siSDOfm73E3XxYrq+FA0pkjsGK5abW9yoa6f2D2WHa34rDstjZO3orbYw
mH5JOIDyY8nERIBWNdIFcjE8tkiH0cMWL++JUxoMFs1YknBtqQALzHVjLmo8g4+Gw07SjVztVgYs
jBjV+XCfkwvFmRjGspJKTXfbIBxtQ4GtJRdHVDgODeIHigzUBFdFY7OkWD6lIVq9x8c1sINf8qXU
ALHZAj1PJLIqClFDMeq9L9mK3gLyF+HQn9+hZlw2aqrGIlBKxlIX6k3tutQjxG45JgKSjBZYfIeW
eTPR8X3LHtTxFMR4sfZN/VSJo0B0Z30/zCG4zbtX60q9xGxFMZvbAvVFDK20NTccZl3FOGiW2Zn1
BcsJD45wasim3v84+jSxgrpcrDT4A0acAVJpq9dtmiZi92ulmvcKIX2PzsWSqzV3wJ+hDeWFSGgv
v84fglDPMuIFIxOa1vb6+YXLyWUEvrakWuRAqTM5y895NllaNixaAJumSHqcD51mbQkuFxfTLYqy
XRjP033jXSK/bGEFkzqYXUTwVCoKasNGPVqgBoQVx3E+2blaahy6cZY0Xk77H9dwnHnMMUUa0NCR
s4epMAwwdNPjscdhJblkclHxCREZTFqHya5UrM230/HW6VU1v1Fadt06uNew9X/3twnLWOJCpebf
tc4UuTCQZ1qOfdvgDHrqNUtEAYvQ9RIhb34xjICEwh4cRDHyP2yoOe7InIxQJlm3DJcL6RJPsPW+
9VBzsdlyUjMKZeGI6tZ6TspW645I5d0KGRSLpXUYQKSRsmJAYDnfLCJfWlb232yx4IzPTMtwixhS
ra4C+dBBuZhf0lamRwkzMBwoUavX6o+J8w2ep0aMVdJvnE5yesHw5a+2qhdxlXTCY0HqG5RB9KfZ
oT+ozb7+q0vVQxNo+hCQTSbNf/22sVW5mbY+/0zrw2T1LmEVTU8UQ62/nCYVPeBqa5Jd4fayuve0
790pPV3O+exx3EDJ7sTnHB+Yg24DyyPdV66DQcyAP/6TGy3aj2xpPo2jhYYw9sPVZ5VQxdJjAhev
OdEIZDnt1nFliJe81CWQ2Lgc5gpgIEkXvSLNBnIL0vqToFfBTxh8QyqarwN9Zlf3KY5PcXzpy7+h
pqqLhmNC4ktElCqgbsM5nLAzhGQsmbHlfnK9nF/HEfCkePuHBSA4RhG93WZypRd0bqxB2/SpAmhw
DE7kpMFdDlrvvmI3se12riLivFbG9mg2WsYNUsDgaUpxSt4HRVsNI6quCBZYGkKwZ0/RODRBxHuf
FTIdM/HpAgmwuNp1jRzJloxswPN9bgQgif/aT5StcL/ppt0QCqymElW95Hxj4HBmuze/h5Aqp7j8
9UmAV5mMuL9WOx3zgyfSj7rj0LMVb2w1fvCYqA10zaI3j5TTvOtlQ9JKDdpI3hWeONjiShAwiVAE
ULOHii1F2wa9ALhARnhcv+nXo+9m4qg2hUk3YcNsirj8Bhu4uPs5VM/c5YneoclxNKoJVKLaAZxz
0RIaH/nXJcTBKauF3hwgmo6uW2JOzLBkOi8UJYTH3uRbtW3rBr3yQ3Z27wqJBFARkxQfdFsgXnhB
mVV+Mk9lHrjILvKDcStQL0ga9kLdkEFPzyxMwDxryZ+pBb5YxsdvIsI4r8aWG9X/B07QExholyKY
rfmgzQ4988UnEEcXouQDkF6xguVuG5ipmoWhmO4jSR0Ue4K0pBFq9HDvTHN88iXY3yzAIx7ObWis
R+9g4n7KZ7m9Dcz13cvBPDcX1uGXGKHL6nsdg4/9vS23ukzrc+vGmW2YtRMPHqQh859N3wN4OylK
rBPV5INN0sp8L3FbsTWHd+hbg1ag0tAPg+BxAgkYsExfR2Kz+DKJduEHL5R1wxOE/HqvdxSlpDvY
r3vAAqgEGPwmoE4iitWOtvG3YAfQPCUmZylUrnYe+WQKHCc8XvPSK1aT/mHKPnoU1xQfr1rYMNiO
2OQMeVf3eVjdHSMY42/OPTgriAIUnzvlvHs6PvjRONAKzETTbBfAgre2IYZU29B5/WGM0CDJ2Lvl
8a2VaT8Cw0aiO3faqn5VXTer0YH4tKcUarqEeI7pyz/fSkEuYjKFNbGup35pEfNT2FMLElG2PPwj
h42oo/4kr+enQM7v2LKL9scCMKCVVbqqBsvwE72ZBiypBxpl0kQW7q3yfy+7tciY09kgaBg9RW4h
XnxivtSTjp6uQ2a0XUo+p4OJltl943wCzE9ctoUwYkZfcczj/5Rh+ZLUW2RtruSKdlGbR011Lbeq
MFkh+uLV3KjBB9rOGuH0v8kHk+CKR2K2K8LCeI1Nm1GXcKNkRuDYA5eBRlSmLvDo1CSVpxSvNpO/
+k/xm6CSTKc0GJpZTSrK23aGRwhbqphpAi9rBO/iAq33O/G3rmo4Y0pZwA9MgbR8ugcH4PvyI5zI
kmxskXyvl2EiTtAJ93C+t+w8axyGcyK+OlMsPp7jkxo22aoJXFMlaISdHL3UzTgVtZc78/53VwWN
Wg3hUMBKh/Ucb4EkFMQ3FaLtjtYYatkkKOj81z83geNik5JFJOUlLPn3hFlQ+XowFAwyvTiWBhpq
TMkc5T0e3SJpWWcNNEJkG1u2rNqWzkN2ksver3pjHYttas+zgj3CZDOOpojGtxKuO3zPtPk9VW1/
BUok/r01HFLYi/aUxRvI2qfqDHjF1uQ+86Tkb/SGjwcIti1iXUYPd0yRKs45MSr1+whFZha/bBeR
xMHta9MTVeZ8dE8w9crTCvAx9e+w1AQ+wGPmTzhwFFOpKLYP89Jjt3fchVPEXZFeJUSkscQKyAnE
Hz2eZ6j9UI05H4yfr75tMgt/Mvw7Sr9m6ZitMC8MpjFbqfqC0h+R8QT1bCikUzQhmgXLNhmOsJ2V
PKkg5lWkF50Xn38dxCueawdSNGOpIg5W7CYKP7+KvBy050AfvJaLz48J+pR5bxM/bqEEkw3otHOr
K7oBBkOLd+0EnpPSq+IoupiOUcgQ23bYe9hNIseIg72dxzJLhnin8tkvVaUAwi5cWyR9zYhHAGYp
sq9NgJH5x1EcZGWJ15RGmeiS3nRy9f9J6tCBzmd0iwlsFKN3KDZdTYrpibxBRbCnrjl3Keq7OvTs
GbFhLjq2Ti9q47Z8qY//WhC1xee5TQ/k+A8Hh1B2ZGgNn2CE6Bpo85juIPKoYC/Lc2ZkUyxagTnU
UTjsSUKoyDKxu+5tl5dDNJSkL34ZKyNFyh3Hjw3BWFTXsVE+RR6eWEzwVOPLGK3rROQpTmNUQcmd
HsrioMxCA1P4hYLx/KjNoj8vjdd1VlWXetz/hjNkDl57/IFk/Sexe9/Omi33mhe0iN9qrWhrpH1I
pTvdA3M8Zaug3cASUU6i8aK1MtczsMDRAII1noYYjjvRWx2JDsDoLhxa2fiTJUxcH5VfKMja5IMW
CnQC6LFcBUJXKlfuw+KsPs9AugY/0ZraLt8Wfjl3xbGcLtVZWqPpJtpcWqrZo6F4fnpbPbzEw7A0
CagVCMHM1daz6YZjeiXRVtFg5ETS6B+an99Pv+W0ji6QK/1PPNT80lW+xIR8Ja7MKiKDJGIUC0uV
ITMavurWGa+Xvc/zPGLa2uvre1u/6GV1cxlxmvaNvlw/EgxGVNLsXbrczmu3XIQ8SEy+el0G6cL+
KNQR14Rgz2cUojUD47KtQUw2s8Fe2HvZypZgbGsFfCEfZvLrIDUJhK2S1wXP5hyO+9lj96tFxF9q
D3bqikN8Ddx7pNlsdHGERMNTjZ5vaE6Fl6ldGcAkgy/ssoAh1uMQLhy/Q+fNa3s3xnYR4tZYa4x2
Cfvxpz1C8jFxeS/vjXsAH4m5xXz4GsM90mF5wgMaGMM03a/+P4Zu74UTGA3jwbpqmCwAoESv+SME
zIwE4u6B9qIDbFw1emEnMiHKNOEX+1PCQ1v49SifD2VK+HMO8hrQgY2yk1y0zk/CVxEwwbxVpl0d
GnYA3kZfOChcr8+a6Ee4qJNOXXYiGJUY6tGEx9zigJ+JPZU+Ma6PZIacPI19fATp81VRM/cXzd8K
UscSd5SAA7RhemfhDX/BSrC+TnT5Cw1pI2FcrP5PDekG2NBW4pzpIilasboxE3Gtpf9P5hJPcrIe
4xNY9oKIHWL8uUw1d6KHHfVACMByfYfHCNR6gnFXzo5zLBZgw6Zfn9mlG+Yg8zEeqhKeeHal12Wk
NhLB0oln7xsN3Hh/3ahqBjUxpwIZx2VcLwKD11qGxilkipme7HF6Xlq8x9DC0TLnnvRqDFs4Oean
Mc7/b0gnd8zU/duCs/a9IPO0kwN2+4U5jFT9dHuRvcfgo4nG5gkGjAp/xYJYbfhRPO9/lrO3OG/e
2Wp8FwWVT55hwax2m8eIPdYWJC8XTlXJ4upmEX3gpqGluOdw/T+385Onpse+eWyrM4UTJxJoRc4x
D5yMKgoyi5GMUY/DWuhqoHMd3EuYH0mBxw7fc92cGftfMuqhKVHDxcNnARStX7A3Au9liI+vrsiq
i3RtcX2tng7qpeRISU4gyxqEF/H1ndjvmMyN9gqp4pjUYX+YVuPgsah2/+7yRW2v7gZr8LJAR6nE
YwmqdRIbo9iWiXlcn4kPJdnRnu8Kc+vVSd0+Qxw02rXly0dBD8eyrx4RFeeoLcNE83BdFb0vED7v
Vh7Ad2Yu2XwAvyZsMYxhJ+BhigV4TBdcl7+AIS8az+4QpmMuX0Q2xEXu3N5Xr/+iq+lDv1nlqEUB
e5qj14aJcUSPF22lQPMtoyO5uCCOOLI3bOnrv374b4+xQuaRe9HpRpeoPhCdRd4LtcdZbF0t8Eal
Vife9kfimxakVcddtMsqin9ZMVZTq4dRmcgtptTbfjMgCpnUqQWzkGeMN112vbhu8+smtPpywnoR
JxDokaBST0I9/OoFnuIp/qY6n7TzhTgc8OrWrFJbsF+jlPLCCI0jFX60WZmTui9KYDW2a3B4Xm1G
CV8rd0W1VkCn5blPLUpGbhFUURQzJ1hgplYae3W1Z+nMUa0ovRQoloXcHETXWs+uV9k/hRlOdsCS
wIEb+Nt3ER07rxB6XZRtFuKEl7jDMlQmgwQ2gDZ7jKjFW1JQ/CeVaZ2pXct+g9E8r+1YdHdpDGkm
aRhK4WMN/BpEI4JBVi8XBSeEVROouxDCHeTbQojhycUDHDFlgMze7u4wXIC8S/ts2jksGU+OfRws
EMFT72lZd49+ZfOcS2qztfDn/fdowXeNt97Y39qe5/cMkttgcHHWpGLjR4X7OWnqWFQJkg/UDEx7
7hQoiMgnYuwZ1Z5OVpUax3UprhzqVdnkH6viBwz90M18ywK1pM9rTGbPix/l6z+i09x/Ju+b9DhB
04ZE+RRU2amduxtm2YYWVCL8eE3Ve+Vf6CDnwZxfOcTCklDiW3HkSofw/rUe2qKeCkZQ5jU8EDxr
B6DmFa6PygQAZbtbkkL5a4d73fIYn9Ehib90qBJUD/4033M76j86Js1ZpIBf8DHf+UiG2XjKeruZ
+kWYlQC52kCi9nvuckcSpJqei6HNfLSYleb0cOYdo+8QY0rkCPAsaULIczWK3CYA0fCNjl1Jf1Dj
hQr0ijcJ5wtL7GHflnRcowNQ2uiKh3xtB4UEGOTF0ioqhG2jDIh9eNdQ6MfHgWvv01lF48n4PsHg
Xhxmhf61VdXWU65tApFooDqvgWnA7fTxUIz1qXVVjoeZxebiXr3IvtIUgtlzyzQLAEXkf9k1hNzM
/4+ZFOZ8iG4GFguS9voaRYEHK7kRHnlplFjKit1n8W1bDTSUQwTfYlGyvtT06cp27xi0jkNkhenH
pD9wU6Rx88xMwXyC9OFILT+84IcM+wHr8Y0cZluNZS4oBVNmnNK5C3p25fx2BsU7+F9ehSf4xyKe
FJvEHB/Otm1/V8f9J+lFQZQgjPsPHOTvcGy9tFtVf3MNgPR3ROzWlZxsFUazfs+WmHJe6IZf9nqA
lxf97SatcqPVfmcBXKrrnYJfxLFZ2/5mMncds1Pnan48H05T4wUoBrowr7LgPPdI2OENewr+81jW
3815AR+xDGxBbRdO+7ZyxUacXBiQducLK9uBovWiwhNzGBYnEdHIdf1BF5p9/cmFV3PmHlTELG9r
dlnyTqjqnuB3hkCsG0SyFq5oGBS6B04vcBYKQq1P9ZPQMtaO/uH598yOqG2pXX3W43Hx0AhG7v5R
npvs1FPrB2aftBK3fFsTjry2w39EPjiflg48dMiIfba4n7HohllwZSiXKt7DaqiaD71xqilk0o/c
spjh4w7AQaUgGM03zFHzGtPkuSpLLU7OHQmAfJV4Hgw+BdBhknLseyJ2FHzckzXvVyWDzprXL1rA
VT/y1P30/Gizll58x8WKaxcR+LanMNnErOUe2JmYR1l9ON3CzDhGMONrJToGwbxkSgnuu8T/Nbzn
ZB5Ih6oiTknI6Tgw3/d0TSH1MIgGMml9EwEOxzvx+EmKsp4w7apkemy4SyrmLeighyqm2nFzaxd4
QxszXblq2WJvGLTC5TyVxzjSNAHD/FmQPoJDGgDbJNMSNG0LKTL/6I2voRY8KypW/aOdDauWa3F1
fDSMBdMQeJ0kwjcj+RdB9JW6jW4r44phSDNpsubZoBitc4Sv2AotKY0XFzY4t1CNnmblhxItqimw
9oQza8fTKR5f1fn0BFCbBMrBD7/rd9oaZtXz9fyBoy6mxOHTW2YEJ+MIBJJxlWRsVyubUtAuJHjy
M8eMLlLhRcBI9hAJQTTXGnfUuzw5b5DdsNf9h5ARuOXgiARmBcsLwZVyVVfYrla0B2IqwzXNcFfR
IrIKSVgqW3NzxVci4AaZ+MIgcYVGYoHpkI95H+yJs2CXoXHE0VO/dZLfnQMAeGIU53EoZyZqqFbo
w4UDmI08v8+QNAqbitAuUrLCMqBNg4+w6LzNnJz/D7IIOLm3seg0CKFx7TzG/2vCbw0bCoRbS1ta
XjU5xaRnwJOmNRqyQ/14rH1npxyuxxhjqDJBSTB5569EAO+ZOyTS3PUpd3l48RG256+z7gLangLY
PALr40gdSBLTuYkUeMkuO5Hxts1jpnKwSdsXpQ+iyFoon8oFnkVou/yZ/OJNNFbWzrJ/aeyvhcVr
41C9RGG7oWZrBep0paqqPOvhVnIh1UnCCP+K8/F1TQWTSY7cS+dHJbxseW9nXLdksC6BimsopTh4
P6VVlWZt0d0fUemh+pfA5Cn40M6B5cD5bKtvm2GpMCDQzUb5Q2XcJH8BgltGsD+IijpHE2j9r9WV
7CYqD8U8lYOnyZmhDpM6MTKDI1NqPysptzTtBtwdAYuFFc5+cvBeVzAmTphsCPRMkG4hmjq4oGSP
G++UjMbuVjKnlGLPwqvwDgZmfe3P7EgOziw5Np0vF8YlZflpMf7cDkvGBpvV7xEjH9lau3Tlm2Bo
b+J41s+40YpwbiPakm40flE9S/AxETuSVt18R/tO2zplnyQsa7ww4FBDHdWR2bwUSenOFwvEv1uS
U2eJ+dN+CgbMo5ewPCR/mL0KHK1bJYNOu3K/rteN6gv7EuazavercZPZ8XTDpfR3zzNJ2AgAKJfl
p03KUtj3RoehCKX6r94em/4WQIMLyqANDiDe1iLs4hiLmgTrPl3fZ/SbPsRcTpOBaf7izRDLQW9G
kZ89lSALmZ2wdNd8XYeoD7p5GkdKqFkhy06gheQRC/SMLOaua/jQL4TDhXikN4xdaChuZTJm4/aT
AFch1JjAsNURLuOJ0vN1F0p6zS0azblw3UfmSSDIpVUfBIgVFxd/OZpcnWWINozgKRgCpBFPHg0N
xR+WsEogFk8NX+9yGSIOORx6hgfiGNLrquKbRGCacJft8FZQibWVxDVj0oZtwY3hJwnnW4t3lgoh
GY/S1Mz2/UeyRmSjjUPOgsHQjTpAxFySWI2M8TxsNhwlHq/lZ/f2n8+bcY3oTsu5Iw+WMRA3maH8
nuQRJlSe+yUMCsUOQUkqIlOGOrRWz6aMdSzbI/4z4mjZjgU9lfn7E3oCVMqfbyI6xr7H1JJ2QdqZ
c0ropHNoWHqgqXewb8kaEM/8kVQBqWZZ2XMkteeP9Xcju0Jttl6Knn1gHXRBbss1hebNzg4QcvCO
dLIH+9hez6SYOqCyTRRpmyYbWyF0FfWZ1F8FrMznf/Tsguf+vuAFjxbshxRI1yvJ1dsuQpfQPJdy
wYUj7ug+KY6B/cuFcRjyzOlXk1yDhada9dz2DDwHdtSEA7HXkzQO6drzntWOAYKJuVkhuxDtoAIA
YOr7endnudIB+x90sgHbadduReJtvNG5yuFVT5nRQzPjk2WD0bdFv43EzEM5CUo2EMUcRdu+LfRo
LHzgsCiMRxfw9XlSph6JXhDOsdEVadeW8LimYrEksdMW7XVGE7UA7AQQoebKFGZFN7WLMsMfXO8p
5RsLzQ7DdVV92c8LjspNS5lG7RW2vDQP+HXvd68fH4w2Q78wWmVqAfnbWO41Vz6Iz+WLA/2sVNyO
OqbewZSCbmOdHLhz1/YkO8CQLtsophvvKVEiA15mtRt9kmsh1O6B5F7ApY4OpT/VQHF/kwMC+jk8
BsBQw5jL5WKSmWxmg//0716JeRC1RKnFFdpbED5eyBkM3z9vKPOPtBk9NgzEWTXiTJ5bMc9MCavq
36Smvr+7q8L0DkMwhDn/fXUMJtYr0PByYk9CAHMBzwDHj0/N9JukcCaIWzMlhFVjEn2Hsp3xh2+7
bO48pxTW2C+LUEXHziGwIAhZ40gr/J1yw+rlllVDGsmJf9DJXmBNNqWv7ZtcW9VuvBSpqcPcvlX1
/SpvMNJIZTBXeMAgKOBgMaR38L+0QtQs9YKs+k7aVXau1MYox+gaZhw+UXc1nVTKE5a+IxMZEaJc
jUHPwcbSlRVxiFm1zKiUgpjM0mByecLMXBeKcD/Wqa2yLU0/61+41hAOTpRHYDNsi9WfURFkeW7u
IClB8hkWvfTlE3aB0JycERGzjx3N2krhWmaVyv2iYC2bSfmZF9jnQqhN1JH4n/MBbWgSmPGdUuRE
esXevGz35lp2E/KbN2aEIjVyY3kknctCHTvDClE0iaG+jvmtBzLKNtJpOs8mQrZSHhE1trVpziR9
k+cdbbVxTO+He/LvzWd48aiOboRPYR6/AAghDUb2Q1k+NYDv0IMxHerTchnuFcgacyucEkHCYlZg
DQ5suQi06jQHeb8Xz7ezmg9aK5I+whTVVWLS1fMzMI9HSb30yGnTrRjSQVxuH/6/qTex6thCf4DK
M6kr2N2OR+GenzWBVJyRKEujiQ2KASMEsH0Rp6qBLTpYCNXTwnyjBY433M+hbI9BCKNLd4ARDs9T
yal2VyS7rYK4n4IUx/xd47ugNsklsci9aBGE130uwzlqJplKtj4u21hpuimIZBVBS/dDYDS46ZrR
SqllXGXWYfHQpszwBkXD8zJUBZkIv7kD6D8xcvmdlCYxHXmbJQxHNavxpv4HrzNGR7BHyGVlZyHb
3YGmxN7o/h3JWKAC9ut74fjRu/G0VJUDuLunAZ7O/skdGiLxGtnqJ6948256a+YXquGW5oRNDZJQ
80EIxVs7lv+JxEKqfPf7yZoV38ZCCuq/sQdtCB9tvPcjQ1UyEtLXgLTqzQ0/Uk4lqJoWS+y1TICz
FZK5g4FvvJqmgZD6jzsbFhJ9PYyJ6vTaCNoChwF1PKzbBcsZzk8JWBqSEaIhmWs53L/tzMRdMDvZ
bLmiMpo5ZM94CD87MIW+klQyTQx4tTgbKDV09F2Gf6e5EVW1zDhmwY+MlzU1HpUoTSeApK+7FYMD
VQs2MpCrhMsipY+IDzH1nMcUx23i9CAtDbD+2jn3V6SYNuYEqbT0yMlqj5chk0Ik1DGP7mnl8uTy
hEIfZNTFBSrWB0KQf1cEpO2BoTAXVwC84pCUD6XCkzvVP0lkzKrXZZZwDZdGLX8Q9DCr5gtEMrdK
1Jn90g2GgR33AwbdSXhzOihzNs4RTKgIjqB2+G0ObVJRq+cYfdus48mh/QAuBax29KwQlqE4KUty
KyX8RcfF5dsT7IdgiM22L9mK0qZcromfs44fcnFtwZuFOo+EzzdKu7jtERboR+aUdlyyt0gd/5o4
KePFYHpwaL0hHD2Pij5Xqlz5F0VTsLB5qxvqA2JiqcXdIXqr9v+9wFCaiiDgSFPANwAcWDNsqIA4
O5RPzS9GjtShMSlgzp36BXTJqeuMAlk3oPz+/wuOa0SEBo21XWD9pFF3JAZH0+BlRFeowcGibOAO
0ca92/lq3t4OMhfEGXnJv5hZP672hbQL5NEpOyYFBCR9CxSEMIWJjjUvtAQSZmW1iTicjjjB+GmB
823l4VBJ7AFGYPSeGw6YeR/m/RAp4uLviSGG0E4jdxSG3Z52PPsxaZK7dgB5AU4lIk72eciIdhSZ
kJbU5qulQsww2O3U6uI7I5aSWQE7ltt3/TnN93xxlJLCmoEWGqIYnY9728610kyjPfvP/VsDwslE
Blw9a3/SYlHaFGdSCfkcYQ2iju2HpchhxIzUfsOT8IB2sguUKlGPcLKb17Rq+p5lJUF4lW8yjwld
s2AeqNHsSZpRb2rqaAq4MtlBY2nCA8vhdJNCyOoxRHgcSfPVVEhIqGVJAUYGwchC2m1zDymdaX2j
fottfpMDOur7k2oQoR4Q5OLBEYMB6q64EIVWiDpihQg9XAuaduSMhZGgPj8tckjaKMMH10Rqaiqs
5jpSsJsx+I8qqNIDtTpMsET1jAae81yeT9adiD0uH8RB+IMJmgyEJ9YU+CfwRHyOkZN2ctQnnlhW
DpKG8NY+P13DS9UthTieIZ93gBnhoqbVNwSdLFhIu8jemBPVNEU34HaGdxPiblPZk3fd7wPSx7M0
oKkNwBsrVSOB9fg/4C7/XJ+Vs9RnabsSOyHKDioFXCQNuLtBIHH/shMGuHR6nuIRIQI99CvIuu0X
54HE5whKaP1Mw5vWcYXkYIcDGmR134MpufFb7kW/Cp+H5a8DGlC7RCUoBoGtmITJ6UkJPExZZ7R2
ncNKy62LFttmdbnJzlMGek0wpZenQ/ALbm8d6HJCngasaaslnqJgObkpvWj0kIOcVZa0QLi11Z+3
C1OaPyU/AkIwC8mnSrh0KabFkQO3+N4lrI6yW7EdfiEBOpuxFzygW9wA8O4MTbhFQF7oCrPHVHrG
JA1+JeShCE4ewvrbccZeJDt6UcWC7MJgc+zFSXLKW0eiwTlJqzJV7gDz3TPYcuKUsrmfBPgtUpLh
ofv2yaTl3EHmV6rXr4CD2UTQH2x/SZDigGyBbEgEn0coMt767Bh8UddrUIm2mc+an76uOSJLbVCh
6j4SbVj9tv+N02+exv/igIZKdeLscET6yc7RWrKiLtyVzn7A8eFAi2bsBO0fzp58NqXlz9mfyEl1
TWzSAV84U7MvgyvlMJa93McrAnIajb//MV+rbWLCmAkfvCKYVIWN+/SSNKIKl71yA0Wc9+eZQYAk
AvYISkIkh9Mxa4VvtkZNrjTtOlphSuM9p2mYKoHtCgbMrecrWwH7xPBTAIyW9elUB6afFob7Et/V
ClZ40m0sbxteSw7fcbglINwGkP1xcKBBNzizIPKH+sx42e02QF/8Cx8Bh5QakxusPlkPBFkB1t4h
zxaZCPu1C0M6LXC3f5bySmUaoD8L546/E4pZxvQI2wdMpXNyZH7dAUMWmHetLGjhD4ydUJbcVk/B
hG9k5FLgunW9/iRiwSKyEmob0bMs2AcuK32r3MxOIlkcT/UceD7Txq/CZPaukV42qcIwiyqBdZ2I
x+HFQM8e48NsjweAMpKoqZHR2UwD+PvHlXAkarVECfSXs11VAA1Zdoj1ySWeAxoLMknigGZ+2iFQ
bE6MP8OYqosPdwexSXg8RItvgmGtaErDN5b5lTBmVlLhTlpltiGrGooYTAPezc4S/CTfM1pRrnp4
t21uGp7BcZ5d1QYuGrm4LDCRf9cbCU4DZsBBwfZo+O1JtHclNfF6d62H4FuOI8fw50DzZHQkqJTF
cPPRfGZk1e3CurgHuXFIALouLT3id5vAH6MVb15BL8vXZvDXdZDc+Eq1ldD2d8fPIjBTorx0I8x9
hvpHfwWlWZUt9SvL0Q2T2TRuhJo6ReAgZzeg/xGAGvWc4vpMQygOG+/IvSoYqwJffXa953Lyx5y+
BNNh1DO17iYEUhSGW+NeYjFIcxviskV42Gn6I+IvdXBFo06E84Cgp21TUB0Ti5a4j7QQRuXG7q74
eVBrpbbRR/FV/WSZN94bpBhEgV1LLwFSrVBtjoDSYgAW4lL6Xk4ZfZ4jZnycKZRHrKGOXqOFOceJ
snmouNmZh9xZGfGnurWo8rUkGrVBweZPeOqR9ZPv+mUlDCBvqvmMwXb33frx7uBFJmDXE3X1gBL+
LVc3dV1+t9W188uKUSHMb7QbjRoUJCEjd4y0zsgY97GkPXG9b0ovTQ6kKW5IkvnRmCZPXHS+qbJy
vVlScFA//v21rODRPIeD7FOHGwiwKYpEhoGoYjKS/cWU84WBu3ftB+Eouk6dIO5nGZEL+zUdVRu4
54i/PLmVaLQpQiJdstciJUPxWTTn+PFdsgIZ+1E/1m6mMiY9k43MmelYh7Njuvd9/FsaBQdafDmQ
0975Sj7PCx+NRk9BHtC5zN+RboFvzas1jWhGuRVbtu1udjGwembLqmweCJTI0uuYnkae04UrhG2L
B8x2R40kH2+pXSFTYe45UcRrFJ5+HclX0oJKXLc7tCaw4RB8lVtLFXf2D7kiPwofsc3qsOu2exKu
gT4Y7gW0sV0aWso0XL3raIX2cy3wgxo5fX6qxp434HoJny6VVBW1xEBmywzhYzW9SAWULNWyJkgc
FeihCjqqR1CO1aYhX0b5wpy+zcWpBscqfb6OnkKPlsvf9dXqVh9h3lRsSMaK/WbouHsNbcEYfdej
KC0e8NOL+x+CmRAIEL61Bwa6CK8VmxPh9aSW6OSP5rWl+muJP5ftYBKp0UKi8jQskwR08oDom1SI
NevLW9FPxq8sFZWTCVUvNko+QRbYjjHN0tB1T9NiQb61keTJc4VjyQjgLcubnVK2UwpAm3S8Bwkq
ZMIeQ8vtsgKC9mPL21QhLcpmWwmSEu7BnQvnHvU08dRHbp7EZaOPmGstO4nkM3jh2ofaZR80K3q6
ahQbjD+LpD5trHN1CVgARxt8CGbQ5xwvrtZNHsaRImLpxDIq+LPl9nyCCTxrKWNeUOLi5mLsHje1
8q1siuP4IrCakPM33HY6caMjVMZDRyZPVLO2NJjBEPurOOvoVLvvDZe42XEsKhrvd/B3/5ZIrHEu
EpapaptQUHQvlA0CvQ7ZlNGki/ioPh8r9Lk1JNYpgriR6AOGEidDVMdgLr9t5nwIaa+IHtduGUHs
2LgKWpp6QuXfAVQMwoYwl/wV+DWjE2nghLHGBTKnjf4ZaUDilvpQpAoYMZJZTREd60ldcInCmRfx
++WTmU3DmB3Gboo6Yk401NpDjOOeG0GjmYnIHXm2ysY2awWtQwzaN1GlNzNiGNhKgR4fppqyOlvn
qYehLM8IK40Qmgc/pCQcKqEaJXp27/iNaXHsP8sjYGiuP4eAvUKerhqko8q5oaaY4NnK5U4MSex4
3Qy0m7kIF3EXrqmdcuGGPf+N+33+UA6npVm+AyshDr2gruY1nJxP3HEqQ7pFhpRuV2jxm73kOliq
L9I6a5pIg9LjuzDWrFLM253JynvAmAvqVw8SJdroxcASKpuPIBgibthEmBf8eg6fw7yjEccE5i9u
eux6+rCAKsJQgRBove8/yK6Z+qbxBPXwjR24K0nf5lOnRvmrqmAeH06fSbTcUPIQGPndpPvoip55
DC4NaxFRDqU8x+dzsAzt3/xsHFN2ks8u0ieKb+mk2skBHCw8tYNTY2knA1baj8MgewSwaXNN4LY8
xMLMa3za8UVUjlzyv/GTZuUKfHAgQKCLZw46jZp+
`protect end_protected
