module cos_sin_table(
input mclk,
input [9:0]addr,
output reg[15:0]dout_cos,
output reg[15:0]dout_sin
);
reg [31:0]dout; 
reg [9:0]addr_d1; 

always @(posedge mclk)
begin
 dout_cos <= addr_d1[9]? -dout[31:16] : dout[31:16];
 dout_sin <= addr_d1[9]? -dout[15:0] : dout[15:0] ;
end


always @(posedge mclk)
begin
addr_d1 <= addr;
case(addr[8:0])
9'd0 : dout <= 32'd1073741824;
9'd1 : dout <= 32'd1073741925;
9'd2 : dout <= 32'd1073676489;
9'd3 : dout <= 32'd1073545518;
9'd4 : dout <= 32'd1073414546;
9'd5 : dout <= 32'd1073218039;
9'd6 : dout <= 32'd1073021531;
9'd7 : dout <= 32'd1072759488;
9'd8 : dout <= 32'd1072431908;
9'd9 : dout <= 32'd1072104328;
9'd10 : dout <= 32'd1071711213;
9'd11 : dout <= 32'd1071318097;
9'd12 : dout <= 32'd1070859445;
9'd13 : dout <= 32'd1070335258;
9'd14 : dout <= 32'd1069811070;
9'd15 : dout <= 32'd1069221346;
9'd16 : dout <= 32'd1068566086;
9'd17 : dout <= 32'd1067910826;
9'd18 : dout <= 32'd1067190030;
9'd19 : dout <= 32'd1066469234;
9'd20 : dout <= 32'd1065682902;
9'd21 : dout <= 32'd1064831033;
9'd22 : dout <= 32'd1063979165;
9'd23 : dout <= 32'd1063061761;
9'd24 : dout <= 32'd1062144356;
9'd25 : dout <= 32'd1061161415;
9'd26 : dout <= 32'd1060112939;
9'd27 : dout <= 32'd1059064462;
9'd28 : dout <= 32'd1057950449;
9'd29 : dout <= 32'd1056770900;
9'd30 : dout <= 32'd1055591351;
9'd31 : dout <= 32'd1054346266;
9'd32 : dout <= 32'd1053101180;
9'd33 : dout <= 32'd1051790559;
9'd34 : dout <= 32'd1050479937;
9'd35 : dout <= 32'd1049103780;
9'd36 : dout <= 32'd1047662086;
9'd37 : dout <= 32'd1046220392;
9'd38 : dout <= 32'd1044713162;
9'd39 : dout <= 32'd1043140395;
9'd40 : dout <= 32'd1041567629;
9'd41 : dout <= 32'd1039929326;
9'd42 : dout <= 32'd1038291024;
9'd43 : dout <= 32'd1036587185;
9'd44 : dout <= 32'd1034883346;
9'd45 : dout <= 32'd1033048435;
9'd46 : dout <= 32'd1031279059;
9'd47 : dout <= 32'd1029378612;
9'd48 : dout <= 32'd1027543700;
9'd49 : dout <= 32'd1025577716;
9'd50 : dout <= 32'd1023611732;
9'd51 : dout <= 32'd1021580212;
9'd52 : dout <= 32'd1019548691;
9'd53 : dout <= 32'd1017451635;
9'd54 : dout <= 32'd1015354578;
9'd55 : dout <= 32'd1013191985;
9'd56 : dout <= 32'd1010963856;
9'd57 : dout <= 32'd1008735726;
9'd58 : dout <= 32'd1006442060;
9'd59 : dout <= 32'd1004148395;
9'd60 : dout <= 32'd1001789193;
9'd61 : dout <= 32'd999429990;
9'd62 : dout <= 32'd997005252;
9'd63 : dout <= 32'd994514977;
9'd64 : dout <= 32'd992024702;
9'd65 : dout <= 32'd989468891;
9'd66 : dout <= 32'd986913079;
9'd67 : dout <= 32'd984291731;
9'd68 : dout <= 32'd981604847;
9'd69 : dout <= 32'd978917963;
9'd70 : dout <= 32'd976231079;
9'd71 : dout <= 32'd973478658;
9'd72 : dout <= 32'd970660701;
9'd73 : dout <= 32'd967842744;
9'd74 : dout <= 32'd964959250;
9'd75 : dout <= 32'd962075756;
9'd76 : dout <= 32'd959126726;
9'd77 : dout <= 32'd956112160;
9'd78 : dout <= 32'd953097593;
9'd79 : dout <= 32'd950083027;
9'd80 : dout <= 32'd946937387;
9'd81 : dout <= 32'd943857284;
9'd82 : dout <= 32'd940711644;
9'd83 : dout <= 32'd937500468;
9'd84 : dout <= 32'd934289292;
9'd85 : dout <= 32'd931012579;
9'd86 : dout <= 32'd927670330;
9'd87 : dout <= 32'd924328081;
9'd88 : dout <= 32'd920985831;
9'd89 : dout <= 32'd917578045;
9'd90 : dout <= 32'd914170259;
9'd91 : dout <= 32'd910696936;
9'd92 : dout <= 32'd907158077;
9'd93 : dout <= 32'd903619218;
9'd94 : dout <= 32'd900014823;
9'd95 : dout <= 32'd896410427;
9'd96 : dout <= 32'd892806030;
9'd97 : dout <= 32'd889136098;
9'd98 : dout <= 32'd885400629;
9'd99 : dout <= 32'd881665160;
9'd100 : dout <= 32'd877864154;
9'd101 : dout <= 32'd874063148;
9'd102 : dout <= 32'd870262142;
9'd103 : dout <= 32'd866330063;
9'd104 : dout <= 32'd862463520;
9'd105 : dout <= 32'd858531441;
9'd106 : dout <= 32'd854533825;
9'd107 : dout <= 32'd850536209;
9'd108 : dout <= 32'd846473056;
9'd109 : dout <= 32'd842409903;
9'd110 : dout <= 32'd838346750;
9'd111 : dout <= 32'd834218060;
9'd112 : dout <= 32'd830023834;
9'd113 : dout <= 32'd825829607;
9'd114 : dout <= 32'd821635381;
9'd115 : dout <= 32'd817375617;
9'd116 : dout <= 32'd813050318;
9'd117 : dout <= 32'd808725018;
9'd118 : dout <= 32'd804399717;
9'd119 : dout <= 32'd800008880;
9'd120 : dout <= 32'd795618043;
9'd121 : dout <= 32'd791161669;
9'd122 : dout <= 32'd786705295;
9'd123 : dout <= 32'd782183384;
9'd124 : dout <= 32'd777661473;
9'd125 : dout <= 32'd773139562;
9'd126 : dout <= 32'd768552114;
9'd127 : dout <= 32'd763899130;
9'd128 : dout <= 32'd759246145;
9'd129 : dout <= 32'd754593160;
9'd130 : dout <= 32'd749874639;
9'd131 : dout <= 32'd745156117;
9'd132 : dout <= 32'd740372058;
9'd133 : dout <= 32'd735587999;
9'd134 : dout <= 32'd730803940;
9'd135 : dout <= 32'd725954344;
9'd136 : dout <= 32'd721104748;
9'd137 : dout <= 32'd716189615;
9'd138 : dout <= 32'd711274482;
9'd139 : dout <= 32'd706359348;
9'd140 : dout <= 32'd701378678;
9'd141 : dout <= 32'd696332472;
9'd142 : dout <= 32'd691351801;
9'd143 : dout <= 32'd686240057;
9'd144 : dout <= 32'd681193849;
9'd145 : dout <= 32'd676082105;
9'd146 : dout <= 32'd670970360;
9'd147 : dout <= 32'd665793078;
9'd148 : dout <= 32'd660615796;
9'd149 : dout <= 32'd655438514;
9'd150 : dout <= 32'd650195695;
9'd151 : dout <= 32'd644952876;
9'd152 : dout <= 32'd639644520;
9'd153 : dout <= 32'd634336163;
9'd154 : dout <= 32'd629027807;
9'd155 : dout <= 32'd623653913;
9'd156 : dout <= 32'd618280019;
9'd157 : dout <= 32'd612906125;
9'd158 : dout <= 32'd607466694;
9'd159 : dout <= 32'd602027263;
9'd160 : dout <= 32'd596522295;
9'd161 : dout <= 32'd591082862;
9'd162 : dout <= 32'd585577893;
9'd163 : dout <= 32'd580007388;
9'd164 : dout <= 32'd574436882;
9'd165 : dout <= 32'd568866376;
9'd166 : dout <= 32'd563295869;
9'd167 : dout <= 32'd557659825;
9'd168 : dout <= 32'd552023781;
9'd169 : dout <= 32'd546387736;
9'd170 : dout <= 32'd540686155;
9'd171 : dout <= 32'd534984574;
9'd172 : dout <= 32'd529282992;
9'd173 : dout <= 32'd523515873;
9'd174 : dout <= 32'd517748754;
9'd175 : dout <= 32'd511981634;
9'd176 : dout <= 32'd506148977;
9'd177 : dout <= 32'd500381857;
9'd178 : dout <= 32'd494483663;
9'd179 : dout <= 32'd488651005;
9'd180 : dout <= 32'd482752811;
9'd181 : dout <= 32'd476854616;
9'd182 : dout <= 32'd470956420;
9'd183 : dout <= 32'd465058224;
9'd184 : dout <= 32'd459094491;
9'd185 : dout <= 32'd453130758;
9'd186 : dout <= 32'd447167024;
9'd187 : dout <= 32'd441137753;
9'd188 : dout <= 32'd435108482;
9'd189 : dout <= 32'd429079211;
9'd190 : dout <= 32'd423049939;
9'd191 : dout <= 32'd417020666;
9'd192 : dout <= 32'd410925857;
9'd193 : dout <= 32'd404831047;
9'd194 : dout <= 32'd398736237;
9'd195 : dout <= 32'd392575890;
9'd196 : dout <= 32'd386481078;
9'd197 : dout <= 32'd380320730;
9'd198 : dout <= 32'd374094845;
9'd199 : dout <= 32'd367934496;
9'd200 : dout <= 32'd361774146;
9'd201 : dout <= 32'd355548260;
9'd202 : dout <= 32'd349322373;
9'd203 : dout <= 32'd343096485;
9'd204 : dout <= 32'd336805061;
9'd205 : dout <= 32'd330579172;
9'd206 : dout <= 32'd324287747;
9'd207 : dout <= 32'd317996321;
9'd208 : dout <= 32'd311704895;
9'd209 : dout <= 32'd305413467;
9'd210 : dout <= 32'd299056504;
9'd211 : dout <= 32'd292765075;
9'd212 : dout <= 32'd286408111;
9'd213 : dout <= 32'd280051145;
9'd214 : dout <= 32'd273694179;
9'd215 : dout <= 32'd267271676;
9'd216 : dout <= 32'd260914709;
9'd217 : dout <= 32'd254492205;
9'd218 : dout <= 32'd248135237;
9'd219 : dout <= 32'd241712732;
9'd220 : dout <= 32'd235290226;
9'd221 : dout <= 32'd228867720;
9'd222 : dout <= 32'd222379677;
9'd223 : dout <= 32'd215957169;
9'd224 : dout <= 32'd209469125;
9'd225 : dout <= 32'd203046616;
9'd226 : dout <= 32'd196558571;
9'd227 : dout <= 32'd190070525;
9'd228 : dout <= 32'd183582479;
9'd229 : dout <= 32'd177094432;
9'd230 : dout <= 32'd170606384;
9'd231 : dout <= 32'd164052800;
9'd232 : dout <= 32'd157564751;
9'd233 : dout <= 32'd151076701;
9'd234 : dout <= 32'd144523115;
9'd235 : dout <= 32'd137969528;
9'd236 : dout <= 32'd131481477;
9'd237 : dout <= 32'd124927889;
9'd238 : dout <= 32'd118374300;
9'd239 : dout <= 32'd111820711;
9'd240 : dout <= 32'd105267121;
9'd241 : dout <= 32'd98713531;
9'd242 : dout <= 32'd92159940;
9'd243 : dout <= 32'd85606348;
9'd244 : dout <= 32'd78987220;
9'd245 : dout <= 32'd72433627;
9'd246 : dout <= 32'd65880033;
9'd247 : dout <= 32'd59260903;
9'd248 : dout <= 32'd52707308;
9'd249 : dout <= 32'd46153713;
9'd250 : dout <= 32'd39534581;
9'd251 : dout <= 32'd32980984;
9'd252 : dout <= 32'd26361851;
9'd253 : dout <= 32'd19808253;
9'd254 : dout <= 32'd13189119;
9'd255 : dout <= 32'd6635520;
9'd256 : dout <= 32'd16384;
9'd257 : dout <= 32'd4288364544;
9'd258 : dout <= 32'd4281810943;
9'd259 : dout <= 32'd4275191805;
9'd260 : dout <= 32'd4268638203;
9'd261 : dout <= 32'd4262019064;
9'd262 : dout <= 32'd4255465461;
9'd263 : dout <= 32'd4248846321;
9'd264 : dout <= 32'd4242292716;
9'd265 : dout <= 32'd4235739111;
9'd266 : dout <= 32'd4229119969;
9'd267 : dout <= 32'd4222566363;
9'd268 : dout <= 32'd4216012756;
9'd269 : dout <= 32'd4209393612;
9'd270 : dout <= 32'd4202840004;
9'd271 : dout <= 32'd4196286395;
9'd272 : dout <= 32'd4189732785;
9'd273 : dout <= 32'd4183179175;
9'd274 : dout <= 32'd4176625564;
9'd275 : dout <= 32'd4170071953;
9'd276 : dout <= 32'd4163518341;
9'd277 : dout <= 32'd4157030264;
9'd278 : dout <= 32'd4150476651;
9'd279 : dout <= 32'd4143923037;
9'd280 : dout <= 32'd4137434959;
9'd281 : dout <= 32'd4130946880;
9'd282 : dout <= 32'd4124393264;
9'd283 : dout <= 32'd4117905184;
9'd284 : dout <= 32'd4111417103;
9'd285 : dout <= 32'd4104929021;
9'd286 : dout <= 32'd4098440939;
9'd287 : dout <= 32'd4091952856;
9'd288 : dout <= 32'd4085530309;
9'd289 : dout <= 32'd4079042225;
9'd290 : dout <= 32'd4072619677;
9'd291 : dout <= 32'd4066131592;
9'd292 : dout <= 32'd4059709042;
9'd293 : dout <= 32'd4053286492;
9'd294 : dout <= 32'd4046863941;
9'd295 : dout <= 32'd4040506925;
9'd296 : dout <= 32'd4034084373;
9'd297 : dout <= 32'd4027727356;
9'd298 : dout <= 32'd4021304803;
9'd299 : dout <= 32'd4014947785;
9'd300 : dout <= 32'd4008590767;
9'd301 : dout <= 32'd4002233747;
9'd302 : dout <= 32'd3995942264;
9'd303 : dout <= 32'd3989585243;
9'd304 : dout <= 32'd3983293759;
9'd305 : dout <= 32'd3977002273;
9'd306 : dout <= 32'd3970710787;
9'd307 : dout <= 32'd3964419300;
9'd308 : dout <= 32'd3958193349;
9'd309 : dout <= 32'd3951901861;
9'd310 : dout <= 32'd3945675909;
9'd311 : dout <= 32'd3939449956;
9'd312 : dout <= 32'd3933224002;
9'd313 : dout <= 32'd3927063584;
9'd314 : dout <= 32'd3920903165;
9'd315 : dout <= 32'd3914677210;
9'd316 : dout <= 32'd3908516790;
9'd317 : dout <= 32'd3902421906;
9'd318 : dout <= 32'd3896261485;
9'd319 : dout <= 32'd3890166599;
9'd320 : dout <= 32'd3884071713;
9'd321 : dout <= 32'd3877976826;
9'd322 : dout <= 32'd3871947475;
9'd323 : dout <= 32'd3865918123;
9'd324 : dout <= 32'd3859888770;
9'd325 : dout <= 32'd3853859417;
9'd326 : dout <= 32'd3847830064;
9'd327 : dout <= 32'd3841866246;
9'd328 : dout <= 32'd3835902427;
9'd329 : dout <= 32'd3829938608;
9'd330 : dout <= 32'd3824040324;
9'd331 : dout <= 32'd3818142040;
9'd332 : dout <= 32'd3812243755;
9'd333 : dout <= 32'd3806345469;
9'd334 : dout <= 32'd3800512719;
9'd335 : dout <= 32'd3794614433;
9'd336 : dout <= 32'd3788847217;
9'd337 : dout <= 32'd3783014466;
9'd338 : dout <= 32'd3777247250;
9'd339 : dout <= 32'd3771480033;
9'd340 : dout <= 32'd3765712816;
9'd341 : dout <= 32'd3760011134;
9'd342 : dout <= 32'd3754309451;
9'd343 : dout <= 32'd3748607768;
9'd344 : dout <= 32'd3742971621;
9'd345 : dout <= 32'd3737335473;
9'd346 : dout <= 32'd3731699325;
9'd347 : dout <= 32'd3726128712;
9'd348 : dout <= 32'd3720558098;
9'd349 : dout <= 32'd3714987484;
9'd350 : dout <= 32'd3709416869;
9'd351 : dout <= 32'd3703911790;
9'd352 : dout <= 32'd3698472247;
9'd353 : dout <= 32'd3692967167;
9'd354 : dout <= 32'd3687527622;
9'd355 : dout <= 32'd3682088077;
9'd356 : dout <= 32'd3676714067;
9'd357 : dout <= 32'd3671340057;
9'd358 : dout <= 32'd3665966047;
9'd359 : dout <= 32'd3660657571;
9'd360 : dout <= 32'd3655349096;
9'd361 : dout <= 32'd3650040620;
9'd362 : dout <= 32'd3644797679;
9'd363 : dout <= 32'd3639554738;
9'd364 : dout <= 32'd3634377332;
9'd365 : dout <= 32'd3629199926;
9'd366 : dout <= 32'd3624022520;
9'd367 : dout <= 32'd3618910649;
9'd368 : dout <= 32'd3613798777;
9'd369 : dout <= 32'd3608752441;
9'd370 : dout <= 32'd3603640569;
9'd371 : dout <= 32'd3598659768;
9'd372 : dout <= 32'd3593613430;
9'd373 : dout <= 32'd3588632628;
9'd374 : dout <= 32'd3583717362;
9'd375 : dout <= 32'd3578802095;
9'd376 : dout <= 32'd3573886828;
9'd377 : dout <= 32'd3569037096;
9'd378 : dout <= 32'd3564187364;
9'd379 : dout <= 32'd3559403167;
9'd380 : dout <= 32'd3554618970;
9'd381 : dout <= 32'd3549834773;
9'd382 : dout <= 32'd3545116111;
9'd383 : dout <= 32'd3540397448;
9'd384 : dout <= 32'd3535744321;
9'd385 : dout <= 32'd3531091194;
9'd386 : dout <= 32'd3526438066;
9'd387 : dout <= 32'd3521850474;
9'd388 : dout <= 32'd3517328417;
9'd389 : dout <= 32'd3512806360;
9'd390 : dout <= 32'd3508284303;
9'd391 : dout <= 32'd3503827781;
9'd392 : dout <= 32'd3499371259;
9'd393 : dout <= 32'd3494980272;
9'd394 : dout <= 32'd3490589285;
9'd395 : dout <= 32'd3486263834;
9'd396 : dout <= 32'd3481938382;
9'd397 : dout <= 32'd3477612929;
9'd398 : dout <= 32'd3473353013;
9'd399 : dout <= 32'd3469158631;
9'd400 : dout <= 32'd3464964250;
9'd401 : dout <= 32'd3460769868;
9'd402 : dout <= 32'd3456641022;
9'd403 : dout <= 32'd3452577711;
9'd404 : dout <= 32'd3448514400;
9'd405 : dout <= 32'd3444451089;
9'd406 : dout <= 32'd3440453313;
9'd407 : dout <= 32'd3436455537;
9'd408 : dout <= 32'd3432523296;
9'd409 : dout <= 32'd3428656591;
9'd410 : dout <= 32'd3424724350;
9'd411 : dout <= 32'd3420923180;
9'd412 : dout <= 32'd3417122010;
9'd413 : dout <= 32'd3413320840;
9'd414 : dout <= 32'd3409585205;
9'd415 : dout <= 32'd3405849570;
9'd416 : dout <= 32'd3402179470;
9'd417 : dout <= 32'd3398574907;
9'd418 : dout <= 32'd3394970343;
9'd419 : dout <= 32'd3391365778;
9'd420 : dout <= 32'd3387826749;
9'd421 : dout <= 32'd3384287720;
9'd422 : dout <= 32'd3380814227;
9'd423 : dout <= 32'd3377406269;
9'd424 : dout <= 32'd3373998311;
9'd425 : dout <= 32'd3370655889;
9'd426 : dout <= 32'd3367313466;
9'd427 : dout <= 32'd3363971043;
9'd428 : dout <= 32'd3360694156;
9'd429 : dout <= 32'd3357482804;
9'd430 : dout <= 32'd3354271452;
9'd431 : dout <= 32'd3351125636;
9'd432 : dout <= 32'd3348045355;
9'd433 : dout <= 32'd3344899539;
9'd434 : dout <= 32'd3341884793;
9'd435 : dout <= 32'd3338870048;
9'd436 : dout <= 32'd3335855302;
9'd437 : dout <= 32'd3332906092;
9'd438 : dout <= 32'd3330022418;
9'd439 : dout <= 32'd3327138744;
9'd440 : dout <= 32'd3324320605;
9'd441 : dout <= 32'd3321502466;
9'd442 : dout <= 32'd3318749863;
9'd443 : dout <= 32'd3316062795;
9'd444 : dout <= 32'd3313375727;
9'd445 : dout <= 32'd3310688659;
9'd446 : dout <= 32'd3308067127;
9'd447 : dout <= 32'd3305511131;
9'd448 : dout <= 32'd3302955134;
9'd449 : dout <= 32'd3300464673;
9'd450 : dout <= 32'd3297974212;
9'd451 : dout <= 32'd3295549286;
9'd452 : dout <= 32'd3293189897;
9'd453 : dout <= 32'd3290830507;
9'd454 : dout <= 32'd3288536652;
9'd455 : dout <= 32'd3286242798;
9'd456 : dout <= 32'd3284014480;
9'd457 : dout <= 32'd3281786161;
9'd458 : dout <= 32'd3279623378;
9'd459 : dout <= 32'd3277526131;
9'd460 : dout <= 32'd3275428883;
9'd461 : dout <= 32'd3273397172;
9'd462 : dout <= 32'd3271365460;
9'd463 : dout <= 32'd3269399284;
9'd464 : dout <= 32'd3267433108;
9'd465 : dout <= 32'd3265598004;
9'd466 : dout <= 32'd3263697363;
9'd467 : dout <= 32'd3261927795;
9'd468 : dout <= 32'd3260092690;
9'd469 : dout <= 32'd3258388657;
9'd470 : dout <= 32'd3256684624;
9'd471 : dout <= 32'd3255046126;
9'd472 : dout <= 32'd3253407629;
9'd473 : dout <= 32'd3251834667;
9'd474 : dout <= 32'd3250261706;
9'd475 : dout <= 32'd3248754280;
9'd476 : dout <= 32'd3247312390;
9'd477 : dout <= 32'd3245870500;
9'd478 : dout <= 32'd3244494145;
9'd479 : dout <= 32'd3243183327;
9'd480 : dout <= 32'd3241872508;
9'd481 : dout <= 32'd3240627226;
9'd482 : dout <= 32'd3239381943;
9'd483 : dout <= 32'd3238202196;
9'd484 : dout <= 32'd3237022449;
9'd485 : dout <= 32'd3235908238;
9'd486 : dout <= 32'd3234859563;
9'd487 : dout <= 32'd3233810887;
9'd488 : dout <= 32'd3232827748;
9'd489 : dout <= 32'd3231910145;
9'd490 : dout <= 32'd3230992541;
9'd491 : dout <= 32'd3230140473;
9'd492 : dout <= 32'd3229288406;
9'd493 : dout <= 32'd3228501874;
9'd494 : dout <= 32'd3227780878;
9'd495 : dout <= 32'd3227059882;
9'd496 : dout <= 32'd3226404422;
9'd497 : dout <= 32'd3225748962;
9'd498 : dout <= 32'd3225159038;
9'd499 : dout <= 32'd3224634650;
9'd500 : dout <= 32'd3224110261;
9'd501 : dout <= 32'd3223651409;
9'd502 : dout <= 32'd3223258093;
9'd503 : dout <= 32'd3222864776;
9'd504 : dout <= 32'd3222536996;
9'd505 : dout <= 32'd3222209216;
9'd506 : dout <= 32'd3221946971;
9'd507 : dout <= 32'd3221750263;
9'd508 : dout <= 32'd3221553554;
9'd509 : dout <= 32'd3221422382;
9'd510 : dout <= 32'd3221291209;
9'd511 : dout <= 32'd3221225573;
default: dout <= 32'd0;
endcase
end

endmodule
