`ifndef DEFINE_VH
`define DEFINE_VH
`define getname(oriName,tmodule_name) \~oriName.tmodule_name
`define module_name SDIO_UART_Top
`endif
