parameter uhs_i_support = 1'b0;
