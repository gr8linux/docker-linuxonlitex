`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
meVIbbX7abLNxkVOwTVCmNj2JODLc3T6ALAMYVthw7uvP5mQTAFGgHdmLLFKlwuFNk04e0ERECWK
wMLjdjcKdqSg/KQclHzwCzfxb92vNr637kbuPQ+zotctEynd1R72RidtX2arc1s2djODLQ0Tkdik
vPl1sinBknYXJ3FXkvm/RNeDNuRT3lH2dJRf+EuzIjECjcBye8F4nSGplNNQ1VO+z2rpMLZabCK6
KtusZI955UTjUUjxelpiXKMDNF1fHsgzi/UcqfE+Xu1FjQtte/9f7i+r6i8W+i4q6gI164/7tclC
MEuJw9NsjZHmgRRdpJ/nNwGLDkc3JVLvR3EErw==

`protect encoding=(enctype="base64", line_length=76, bytes=233408)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
RxK1nnhjgcXpw0MIUOysEzN9XG00W9xaj7lF0kuKxbxBwhWW0Npvnqi7WGhwVxTTamIEjejJz7I/
hjvxuJ3w+l1hmHesuVrZe0kFVlHtdxsbqr01S8xVRoA0bJkdLLSsij638Qn6/fFpTMt58eN6fKv1
Xg/6UYN+kIfVBSpNxl5fuuVDI3ZFCjiI4DRMQpCWiTTkaCnqE/+oUPVaGv1EN/YjtLk8t0DLB1ZU
joYNoqiwzpbd/uQTMwj6CoMueAy0wWvSdnjFKWAc8CzwHTv6Z0gdVAZdGsORLNbSiRn4JTLg0BEd
tQp66imErg8gs+hYaVeVFUnOhnrdz8zdu78/8GrjhSpNvOzt0NTqX7pIAgqnQPJT3VUNuGquZWDX
NMY7VIS7Y6619Kn1jKAynYfgZQ3VWnCUeIRmCgfd5VBugTaOw8rZIhc8yXjMM0Cdi80BPpf90DWj
dQZlvcgvbhvXmW/ROyP4sP3yLz9M0sDIrjPssMRi7B4L2lT9rOvlr0FvZyK9NaCEpv7LQ35w4HwB
mxBfvsKcNnNcmzje7F/xLnTy+lagmrJTs6p06KFFAD5P0PI7GAY0GS3yfi5M4gCx4yUto5Nd60d1
t6MtaFaby9dUWg7s+vEUTW1W7UFCLS87+7W5JOrRXmrcWGwPuVSvScK8LwFMF60S4nLKbz+okMZ6
X1+Yb+hibrTJTHzqjyLasakJe3AAXLZRMpYhLFZpznDrvCYmxfWhaRgOQ0cAYTPbngmMqnW2fJIl
+m6V0XwFNcWtJoxtvHd3Tua+myGaAqmLBZSjpncCiZvCTeUzysLeLlWpIQsP+3syBOJAKyUMlsZt
vNhVt2lTWuU2xFAK3gMIiyqGLqJUdEivjrjNIDdRuVRZwXZVxLlKFu1xGgZMB0dsJfoL4PY/skvY
X0o9k2WUhIM8M2lSW5wu2YVV8lvv197uUzyjJf+Pa3tOd6sksijkCFMrdkyIxPOP/T/MuBPVv12A
nUOWy22sBuenK4BfKEgZfc9Tvxb2NmOj70NM24ySgDITmDXmu7MMCVEFEOcH9mQm88yN+V1/TTUK
0ocaf5sIaua+BuVQoXxjYHaOsYP5C8yJ8T4fjXQ9ZhWKnvASwZlruGqliDdQwLeNzaSxg+lyKjvy
orTPI8qFM43xBi4QinNW45nonZ1miTUtJr/BoiVtGtA0nFWv5zYol/rld/vkYSz2NjN3ykH4MDeO
izFTLc73+5b26aV/4fa+qKTl3Ft+olgyNQhz2C1h8xGOH/aY6uClREs1JfMrhS0UNsHrYNmPHayF
aacOIuFjsG2ZHldUp1pq/GVfNjo5dAvDFV5FmlpOHJ2/rUwSpD+4KmcrSeqTTiCNUzM4ohBFT4uH
+8zpyA94yVtwxQwSUAz7nBkHFsF7oYCNQ4AZYdCXekGr8wBa7DcSKBBntztoh3nnbZmZ1+IqVuYj
o2h1Ppf5PcG2vxOrP7iGn8jLmtmMRDef2lW63tkL5Wv/Jm3kTgJr4tDvEE/ThbBYBlPb6GXq82cr
A5MrQXmrohroIyBtxUn8Asfvb3cTD7SllZ/oO1P3ufFP5o9odLS0PvK2RXafhw2W4bBIewjgL7Cj
wTeu+cQUHyJrg36fMa4PDXBy3jyjc+34kLMCvL4RGIexU3j8hSn5BWtpriPcbh3XniAio9olqfaP
YkhNfng3EMHecD2qTsOdRu/8cRJdE1Tftp22Y2m7a9ApuFr45GBqc5BU1gC+MGC8PZBdequqEev+
jwuI267S3OhL+zRbRDQjQmirxd+1HMGQ2EX/qHdG3VOYwH/pE9uxRJ1M4obxeIX+soiFJSjzrhzQ
oL1y8Ib3Z7vHYZWq2eCNAuR04AF6xAA4RfPCjSeRL7P0YF6FQJr2nayWlih2a3nHqWzY89gZ1aTD
Y0TUPH7WZ6Ih+gckL08gz1M5gFGA3ftOn6sw5HX45rJrHOKwL2TIFIAeXGAkCFGgFIen69J7FPbf
4dBNviP6Ikjq6JnPfT1AwQvRLHIUYikBq3bWIpozaSwaIr6UUH8lpTuqEnu/gOl+JpLv7SFt9T05
gTKD36D4/Nn5wasAc+WOUy+x0ihDl8SHZainSsAGV7noUSPQyQ34/WQ0yxx40wjK4PnUyeuAhrMC
5DVDW0ppngBsMD5tNuFVHmOKq425fFKx3roClP9A5cuNAU1na0p9fl8z8cV5/k+m4Mja8ByxzEvh
VrX2QNdm1uF49H2AXhTKL10W/3JpZjnvWaL7ocE6E1KkiCabQdtYM4wAL1m1D0++NJHFQ9YYkGuo
BQ3/F2+qCi1WiWQNWHHI6I/UEnUoylBnxKw5y4r0f52cFvL61W03LnpDhCChEw7u6zwwQ/muEKcX
oyJrvGlbuKiv3k0Rgc/XKcajgV+pcxbjFkaSkNhkReMe1n+GPU5XaIdfDK75/RTsjfr9F6oRM0UV
V+KN9SVtykYMoCPBAJcR7sJmwlTaSlSc83omC5pqBvjxEdXf/ghAaFzICqdYjAHObLNX2XmcSsnX
YVDcvXURZNc/S6/NTWpLvom3zLVub8oJCQs1Wo6c9YwoWym4kAKvNYINuBJgkmUEWr61gjFXhofO
9jITn4v38HU6gHjDzwwYLP8f1I9+sfFhdJfSwJe8r0ZfwB5KZvmtbNNWNdV52wPNJVvKtTX8IImu
FXVaRM+YuRQEHtSY2maSBK1JRU8hGj4YnLS3wzDiTNfHIkxztP9EM7oWYjtRM7/tujVhBfzRx3oZ
KiqKLGQBRXViZ2O/MYAgrZqHtlwy69UB1uZWfSAtrFNuNBRTs3ZkNC4C3ho+irpd2gDXaH7qmf+M
gQIyK1Cjkak6YrfvPhHvnRIv0AbcczEBcZNe8nqIqo5IY88QwOv8BpVEPzsUxqNHIFOMKdcNr6zF
C/iJ5VE036DlIpO89SvVR/gatoZIYtuE2EW7xXsQ3pr1rH7i2NtI0i9wViVMEuLLs9az/0J+H7Kq
YfitvrGRHprrUcgqHBJWQFU1/fTV4ZDa8fl3HE8KUKpOdeX5Nt1r5tlzjcagCvkp1TIRpjns2sDr
9zSjGl7UcZG5O7vZFAooSc8P1F3fTWXHLgDIlhBswTFV0359G7k6a+GdtHNt08Wx4H0OyI7+J2dL
oKLNsTDa1exW/3NYXBQqmdZbhPovXO2AWNDdR+ZBs7nQAlsp8mxbqXxyaMavuhaY63D9F4bgj8V9
6CyLr0E9gKPRUXD0MTzsPQXemRTiH2mrhTgYXZY7frGR34plSzDBcKc3xtohZb3nZcun1QgIaiN0
iRcZwG9miAKRmiOc4tbOQ8DPVflx5nnpvgJqUM00wl/GcSnDZNgpDqhdaJrVhBODstCCzrxZh8r5
JbfswZ8BKpX09e1K8Vqw7oGnrqFLXRc2WoSDauvSuBy9EHEQz5FFMtq4UbvfXjMFD6VnGptKAxCa
a38V7dyKgg9fRKfiS8eS6h8VzmzWivKSV743yE9sB7W8TQXBhYCpwlEmVP59iBjq/mNzFUkOV47k
vgI1PwKKWEGr/P8Iux1nrzqffqje7nPGlWeNrKGNVB29Wo/p6hUUMoFhUpkV/SiSmJeow2jFpwkB
KNuLujG5NFbDD1MrY90LmoUnnf7S79EuLIecPpxOdfKUtei168Hnetg7RsH/CN7d3QuJXX4uI66d
4BWTlofnvna2vkFeuw1ZgPYjv2Vi5uKO7cxV4nIcR2qehT+eq7UDDMSPZ7vM06avIB0RMYawIpAJ
UvCi7tKcf5I+QkE4d1UZs/LJ3NX1s8zKpBs+sSwDApGE0qKfc9IbOirR/Ri+UwVbci2m7NiLyI2y
5m9GcciGn3VeICj8LNNCTzP/ibDHYFIaojTiZsW8pNI8KnjrVpgWOzPUUsJ41w01rgRtkyepn4lE
LUz26ct0zongUDiD7a/xeajvoURZiyFyN7ym1TliaHuH4ujN5jGhMyChYxLYE5nLGyuyMgUA45tb
4YCdPK3xIZ/9DBd+lA6m6PbZ1X2IT0poHGahNmzGHPNzs+giToHwZifrzwL+FpOap8rHMC7PzzE2
6FIh60QUId4x84tJv/mZqeKVD7w1ccH4CKQ0ZaBsE5fmKwcnX16HerKxFNeedzeXc3yWrjXsJgvR
wby5Vr3aL/zhf/7BGbBc/1cNbhnXZXfxlwZjFACHSjPPFBFm5aoWIFjjPjDh8dt+bgjyY/ZtepDk
3n7Bcyk4gnzjywTMSae435jB75wC9bkBBcRPmhF3KIYv4sOE0Itlm8dLHKzUfSQ1FyY5r+/kZp2l
hdzCbAE+chmdUAfL+TK5ZYVXDCQXoqNGOj08DZALAlSi1R0s25yRJ7vv9ihxfT576sFqDAlIrjfQ
h6LXKQkE98qBtXZEPVZWKUJgKemDqZzOm39BVpekT+4ancm2ijgRUQqtgVrK1q1v4DIY8weaFsfd
OoXVJvdnW8RdWcRJashckaEoLcA05oWo9iuyYLrSru3eRdlyokCMO6f2WXJonc/s58L+w5T7qP6n
2w5Z4dWOZVkf99+eWi+V0/qOe795DgsC98ZowkdXzOUWDRudfbyaFLEzJs3Z/3mEtc47waPWSztY
vqjB6dIuTo+mkTL8Q0ssSDOG/uTV3lzdxjxjB0LOZMsPfNC2IJbZYfu931yVL0bEBY8m7idna3jo
0YNqOC3wTJxoz4w2WwR8kiEiBNOvorIYQDJSk8C3K+BxXzzkGb5iGXAfp9bUywp2dwJrIG4nn5Sa
ITIyT+Hdr8D7NRgRkPYRhhqGyn1C8hfUoj9nxwC1izUqQr1YdoKRqmtxREbjsUkNdcMrn+222I+3
rRxehmR7iAnxbzR3aHVlxM0opBm48IvtugbRA+pxF+agiP9DBDCB4CwE7wk1StBf9pSBn3ZYddCZ
tLmEXqtgMvsRSja+nsaB9DHIAKLtYQrlWaq6/asxwaFT5Qfm9NJOuguhLNftxuQNVRyemfztw8Lz
KEOKUZCtEdcHArwITPmKz1o2OruwUpKsFXObtbbygQHW9x5y9W5W/wIqqB2Ns2xnT0wBZeJmaJcA
yUR5Ed++lGt2VTVxjBUDQvy/lyvPEUla+88z1qJY3slz3hH91f2QIXoNouvlam5dqPZ2acvU/Cqt
fdoBUKNFOuvmBnmDK7VnBCL/Shr4ZrTGF+y4WvlWzbUjHhRHrNFg8cb6sRZcSTkyhzCRZKX9nbU0
yycECaOT+m2baRSQwR36ECKtjZe0O5uQQSNg5FqagdwUOnWvdBhdIPxDN6smlZhwj4n7UokKgMM2
h/C05j/26ZDD9KvVRdnVlpm7RutyDG8UqkKfe/0J0gOEllv+ZehPRb+eXdurCP4OA5ugAzLnwN2s
+JdsSedcSoiO4rJZqW6EWV+q3OxZEOHF4lPacWW634al69do1EDlosg7c9CwdEfkKCdQUYqj5eJ5
DPp9WoZys4JbL4VpnqxC6nglUdlxNLMW/C5fle0TEYGynvX8qEMc2srvk6t7AuvOX0bVdjzBZDsN
1s/s8jytaThxKfFATgTkvYLNV5CVxseIYgliyKigfEYOrq2tfSKnKXcQM4XcbYx+/8hGUF6pMfki
mapEx+ad+lfodU4HgSHhK4FNE6mqeETtaAXnALSCZAH8huBVfOvpWXQL7gi2Tmh2/XIrht/+BeGQ
EpYToSDVRzrboRsJwIeZDyNhC9TbjA5R5xOCvTKuRzpxA7YmPoTBs1jnJcMx5ZfF+fReK7GlpOCI
kqR3lQh5lsAKNx4YeEvauQT6UPaSWSquLNl5R06uxTopb68irgLLxQy4a5MChvGQjEA4JyWAX+/G
TjX3IQh6+whgwXcCRrrz8gqbACD+rDm9KwRXJAOjCbWJGYEcR9rVjgnFeYiwgakK68Jnwoc4GueK
fJn9sRYmGw9QxUU4zqaywflcyb68XNU2QJnaEINyHBGdYKU33aCCeWtCH6Bro6ksrEzxxlhbhrTT
8NUA8xUTlyY1KehWP1lWGnSYLS2qUU95BKSjKbIKpHg2ymQQgpSEOIMOfnPYYSUNCw6y+zgPWFGh
vsHghYzQPQB/NITGuqu9JuvzVB8gL8rKUs969vRUO/Y265Ue3GR6CKT59a/4qNekWxb2OiJj1dF/
Y1C40anAq5ST1WL4AtrW5ahU+S7kDBSsD6KJ06r24m2LjfR0cfndm71+G4nNaY3rCMG9k9Sja6fu
ZQCUCtRUYCBqlfJcM4j70mPtyqL33edJIKOXkPoEIbY0qzSg014L2m42RJH9vxoyBfiD0vDf0Irf
J0sglu5fAmqTRKv4eS9QeKS6ORb3uRQh/9ZEM0FUxY1FBYG56OlqH1OgJ2v74HsZWlImoig+QXdI
KkxMSrhkDs1dyjro7CjCcEek6QtlDwZKi16Jg31MSxdgURoE8vUsUc+K9G66Z9Gyqlqg+p0TPeTP
EIxGF7/krBKxCwfyevAybA6geNcYCUnHg9vbvlibrmKoCIZRwOk58fLWN+qMpbPuKFnBPbpC2fm3
5AwHrA/unEuZBximZgzLev393cEoVR1oS5bu2liAFwHWqaRz3YLcfZFlZz1iPh5PDcgZLOf4qNF8
TjL0S0qChYnYwToDphGaPPa4Q2mN07d1QBF6xVdDRiYNz+kAyXXWU/USFbO2vK5V1lo68mTMgRoU
S4tzU+CUoP3Hb4x5ir9yP0xcz+Xkq6kLjWwnK6vYlPilzq3ssx+WzIymgMA0fRsOa8+Dh2TikKNR
Mh393J+vKz8kcmReY0idXuiPLtTvK3Bd++MblGWlyfSzY8VQ5CeeopZSV5nn5UTCSOlFqhvA5p6x
InKpmajEY0djJm55bTOooRyLg1p1ITuu18ei9XCQgmxPiLttM25RAgbgcN6gIBhs4U5dTSTACA0w
ZK6o+lyDLkkEUi6gpW2t1utWCxOEdWsApkxOF+e24YCo+ZYQRdl2aSeYRUwFHVmiO01WE/Dur/By
ZJz+ayxnHiZqSHH+31vehHzk7WJtDtx03bSQGHg8H/cpBVDCU+ZbCIfToEq6I6kjVabkgXT6TVcS
bMLbH8DNkeyMX4p4sJM6nKtEpm+U1wiKzpsskxK8xzBHHhNhaXxM8jDV3awLjmLwCO6avM//4ePQ
F7fjHrpJ/bjaJkQ887q2A3jHrneyxW21u/NecK7F9uZ7duUVHoxetkimdQ4muJbTpNmlezA8OKo5
SkusE7QWYbdeOrjaa8V4fjDYiUJiOPd0kSSDmmJL4VCc9RHFDFh0wRHArvMaffxYyc8hXoWA9keH
iWlweTA2b8HoWIY0D9pTj2NHhjwO4ZYETjBu5RHYiTVsbx3qervB825G1h2H41lPZiOrmHNoG4VO
qjej0D0tgG++x8IDF7xg6idhD7D9z+/AYezgmrto/edqqJ0HOmbazAsSzTY87rqEnNqm5HAuz/rp
+boNze5b3cAkjII1v8WseSEGciakjZ2SqEiEocZfiW3Tyn0xoOoqoYX3whw4tyTy1WSRldC/rJBi
5qstPJmeKscUobSTjcJCqYewCpFmdUpXDV49j+JFIFzkazwVrY8fCLXaUpVSnOjAqMeevRjO4myi
vd+sq56caI7SAafpdVjKc9ckDk1po/NmUFWjoNB5oPXuwE4GzfL1LoBip7XKQX/JYtCXnsOU5vT+
lQrd7m0j6nSQHBlDXpr6KETqdAgK4GTk7hox+BNZGCKKwRb0svu2JREfXPz9sM1nqLVnmiV8QAeK
1Z25JZ6xecKLb0NI665Out2bUFD/X/1M+iOWyP6aBW5WhEHC1TxplGn1vgoY+N7nv2XFkh3/AuWy
o7gYlYQQY4/rLLezgow6Yp0t+RomJEVI8BeuPHtLWwJMVjRzCvmqURcuP++EY4nqKNwmmxiK0meQ
ToF2msDVaUS5LNPRxy+U3BNhtWoRf8eQUSd65+tQwDGYyCX2qIHVXQ7oJ4rDp+dE5t3jrZuhgr/X
/A2BNPluKK8GbY0XMfqScRD67coLEQBPs9z6jrC4NQHGql6a3JXEbNVCY4eBLsA4gzuEKyJ1LbnJ
jwJX/+6UvTDmDmsvnJsA989+4tj1jsFV4ML4vuk9KGRR3XGltRx5M0YRK4rmCncGQSmmtnYFOAKK
Z7IyqwU4pke42kdHc2CTCNE7ucrM7Gr7t+6wxbIjzw6q3aVyPxZvrpyYO2pgYEq9H7+Kx41Gq89k
rwKe3jcKQMwzau9XocxoCZ4wKkWZg2V2a8y+hgNlrZ76CASLV2Y1s01AWFll9AR+yhaRjC9MfRWx
L2HGCfjIfBFKw6X3m/jFkKZAh1alVZl5C3OOAu6Ez/i6rOnIrXihdqTiZL0xkDajLILAYMbmhEx+
Ra4f5iHQiWUSomL3WmqBqGse0/gwB79u2ZN5FQsT5q/RmB9la20RMWWP89xWBymMsE8BsmMY1Pfb
x/C6pmVZIL6WjzxT1Od4g36x8U0XzIjVQhXJr88COpNdHniJeVv3eDJ2xyAGuIdvdQUOwhFkyJNo
8MgrQMJ2hMeErRjhnln/gpWJ2TwtQtZ9QL4g1f9KTkbk3HE2CGEZGV0uhM+zJjuxqu51cnsC+TES
fTraCWc4c/NangCyP8L7zolD3Fv60sOMDo5r5dVF/OIMSVPhLGgUkcNUNE0S565UKmP/OCIetcTq
SWwpwk1i9brh3CS8ULcy4SQMhFctDFLwDgdoVWF2JIh//vXuAxj7SBlwkd4vUYvZTt0kYEmreDIB
ldq4BtBdRUWFI553/2ubvk46jA4HX84mE+/NsL7yVozl661FM5rV+QIKSRemc8M+bVUFbU3dz/2d
BHM+j5Ls6aTlac+2XaFvc3CfrrM+lTtAWPCbULdeKuXnJCTQSt0Fkn3zxI37yf451S5O2YnmEXgo
w9FHbeG7TZ284XJwwADxOYmKCWNTF6Udg3/VvCIU3C85eccM1KUDYOgTD6atykK4nVsS8QKXe4SJ
oB5Ohrrcq9POJ19foWQV2OXrpPZi39aWAR2njsxLyrcEmsCgrCwPZPNqo8L4iaX7expvl3wNJ62X
wqqAtS10FtR3+YdFnFygTKx/UnxH5ImkhWOz2VGA/Fk2Vg3e0myDoCCBpvw6vACH/2lJvSVenePi
yzd8K98IzbqCxlp9remI1GnXdagAULTDA13NFZKAAx+Z2D0lT1KWZ5g0IHH3r77LVZhJ0m/68KGh
rPoGYAu5h3wah1f/0GqsYHhYR2YHMSiJu6agGJ0P3C8LP8yadlKCWhcaT+o495j1GtRNoYO6+qbO
B4UFRy4g47rjwlHyKwJH9uBVGMhpPKeeQ7JnTAW7wULV2Mmn0sJOXwiiWqX86QpGTXfyOWEH8X1z
9bMBFbB26BvDOCLAnOatB2/p2KBxlSFCw1eHxfOxhJW4YYTATEqKckAbrpuNsQ2c2qpnjuSEA99o
M7h9wOfedqr8w6DW21fPyGXzJHv+qm2UGfQPrM4bVucn4i5vU+peTlyJSnT4m8kg7Gw2zIsLK6gk
8ZT9rH9ubW9m5ABnPZdhP3a5hHtHRTwmBp83Ja+chwSJf9NUG+RAmgFK4UfyY6F6d9z1tq3CI55e
dJTS1iW3EdUlryQin5BigRIfeO32iZbUnAkmQDQTUqyt/0tZAFRfkM8HZcoB6X6cPrXC0NDsQv9w
iIMZD7H8Ih5QLCU37tcc+vOUVICGq+eF81l/RiU012kQuJjXQF9Y8Eb6GXiaEcriKS8/LWiWX9fp
ecYeZfJzohB5iJASysIk9gLEn4B5wiYuVJKcxZ0HKTTY3qSI4mpJPgdvRky3rgKwdINON38WcrVm
4K/gsZLbz0FaycHNfzEyDCL3VFUYwyPqDSBM4pxkQg4tAgaF8SEt/4Qq7b+ZsrZxt6LJtyIwOIAb
oicEf0wzPHieASMfeqzhnQApGa+eNqo3DLkrd65JsF2gMCxgFl5e7c7ozZdGNcD1CCZwm3OHlf7M
rNcWZEZrf+4FStYUey2HH1tRYTqlXg9WGnfslU8jY49smvcmKXhdITbXt4XE+5TTqQaIk9roeYy8
faVuzlgawtIJETjUwjhA7FoO6dGGt/Co2np0vIq3R3sexBoIbruCortnijPloIRKCkFTViUuT8pj
h31L9L+wuV7/FzArDFNcSX/g5BmJkCDz0KWC1bWTOpBhbu5RbzzNJTlCVf4ZOcRR05pDNIRD8Jyl
B1QKfKKhteVFzXZZkKHjZBNWBWcRNp2JJtupI1R5gKjGb8Qyf6NP/9U+2AmdaXKrUBTHMjazL/+z
gsEzH4NQjFNgnfwNylB8pFpGfTXjUgK5JTdXxjEIm7ApgYU4ALA1oDiA8SRIHgqWMnPq4wKEtm5D
mZZWnuXVqRqTOxxChmmRkFZkCwm+KIc8UXH5P1xHRzRVpMuz16R5zUGhOakLcSrhvAXM5Bdb/EMt
DXRH2PMali/LBhix8MtCPiSznZ7ZDLrsQjxuKvf6TD6H4hM82oMqecY7HDlMwsWcL2BAb0nqblBy
mLo7rH4Wa8KxCJ5SsoHCNQ3JHvc+9ATSneh6MoQKGYMZGpa1t61FU5lehtxcvl84BuXSVKq3iF1s
F9xkCLl7SCXiaqpy/QROX4P16LkXVSVkH+Nrpx/QUXjT0CWyxlqTlvaCjl22kiko2KWXzrILX1Ef
92Yyq7Gt0ddPM/cBznwnUuqDZcFEE85c9wAfqg1aOioAA0PTs6Tt8AfDvQLVK0yLRxERLORsEM4Z
Kgkp0odz/ULolhgx0jDL0r0gcM/ndZg6gjSl3fezjPEyx+/HGB/ysORtPy8zt2arCzxeBa5H3PaL
YqSS94SpD5jVgs0zGd4kWruapXAX5qcq4mc097bWl4RkIIgm/9hJPINk5SLVUMKEZdFH4L/YTneg
uyQlUMiKByLSyQ/oJA8dw4oUw9Ogip6mf9BpVBzppc3j4s/uqr+m5FB+G72y4kq7lNgp38uAg8oA
2iOVCoJnek4aT6iHXWYdrYDrKzNCIMAMgMqQQeBO26Vs7pyU9jWnWHRORV4oUaWT01SxSj8QVfpD
quRFeno3b1BxAG+xfoi3+n9vhevJJQY857PnyYKOA9/jWyK7WjOQ2nWRoAHvZh1FFSvbsI71UZNJ
j9K93cE66XAb6pY3UJo9TWm28w2zfyf0PzjLaVmyhOJh6lJ4VTMLls22P51CicXycrriquJE7EVz
+g3mT9kC0/FwzNknF+d9gTtJ0h0d/kDbieB12thhNB6ZLbJgbOVLyl1kYkEG0d0+y2PSZVlb7+eX
0p40zCUvcBc7R/QDlba9uHY4eHYVvoD/dNsy2fBkAXXDNOYN7WXVcj0hny77DaPW50yfLyGuFuSX
FWMcvJzNWsT1g9xqQpdEDHLDYAIuMdMKv42Ew7bGXnFUXsYjSOZbFqfIJ+ti6KEmK0+RrPxWXstv
+/13wCOGCUtj+/S5ZN/B5Xf4x6cw6uaRgB6URrvlLgaysWQ7+VgnzUYR0pywBhdMSGjWoPm3HG5t
8DVqrPv/N9pQm9yAaTSICDde7vQRicb6g+Gf6+pgZJMJuMBkzCA2CRzA9Sw9qvNj20ynZ/AEBZl9
t8aWyapaACTXEwr2ef7RYSK9Zpak6V6qKbTdPacfj55ZVKRQUS5vuk/8bFMWHQr0jyq1A1UnOPdS
g+zZ+iEjLGH18xgfbcER1OvdayBRzk8oP+3HqI1qTVL5bIKShT5M/F/axr6WzENnACK8Zw33TZCi
8Qx6ENxjgbRkQtcQ6gRt4+RGN+xs4qjeB2+J4J2QkiAL08onhk4mekq1vdKo4d3LIQ8/uvEq+atf
YynjX6j4sHvBsMZALg4+RgSGzQwanLaP+TR59VQstfy4GjG9scOcXjvehoX9RjppQZ5ZfJvoXzau
i8i4yptUCFbj3lJIkO37z62wsOMgTsR9GxWtE1doNvWf43NbdFqsUq/iblXUiDUrZqNKyWWtR62h
PwkVhZb7M35yQLTWv1+h2PdJ7BazfEaol5vL2YfYmYONwbCx8eeU2MnOKAilYl/x1guwk8FtOPmO
QZCBZFC8mhY/fkEv3fIW0cyP+hZb6Vx5MdpghnFZv7Y6Zh38jslQrRn+vQV9a6DGONQAa58F3ex/
AzGgSe5fUXZ5b6XN5oW1M54m3zbvFM1Vat4B9RgcMdLRaVqeMukCGQL7yWkviKsmhbM3X2V8Q3n4
SBDgZWej6AG2N89abjgHUmLlFn0YYG6GVrwnRx54RJBprApd3KMSGLNVreV1OQ6+lhGR/cIVf8rq
D2wQ98lEiPYhC+2lAIVPBZ8w9wFEnkjoJkmL4KbMIOkUHFvEoA9pEAXT6Nsy7QIQsZdb8G3D5C6y
06NtPQnRuMh5pBHfeTlJX5NHgeSe3Cf24qXZzb0/XJsP7LzsGd+D4arh4FlheSAqfzk7RlepwAqY
aVlK0fAiA4RAIwdy0cBv0bWtJtRtVqlCg1ldLHrsyfqFpg9KxdmfEN8HmCkV8KhRZSfbve86S7T9
LPURXmULN/JleaPBUSgK24zIAxdscH95zLCWUHGNuPQLRg4iBq3g76eVGLTduoFDMQqEu1OFtsIF
QbBwnd4DtVfkebJEhJcD4T6YrJpqzDw9yM2VgT4dp8/XDdMQX1tQptY+qDISXjVkcDrQ9Kd9DhFF
8+C4iVa1fVymp9jIIwZws+6/FM9Hwnhjh3xI6jC3qYb42o1WSdjRp5+k9FKSLDNjaEjDcTr8yMad
YGGWHYoaSSJRBwFG+fHAIVxfpqp4GsdKKebC7DKx8/gsxAUQYHzNdyG76+rlTEDPGUYeRIIDFiYg
LMpdtKnV9kNzbQGvnPDUmoObj18nUJg88YFsViQta5McTahlOlGVrAS8nBY/WBq4/Kkc0zA0Z9Cu
7gBmhQcvPzUoqmbq4wGwR8S1KGNIcTeRio0eoFQzRDVZYDqef/CJduvDfI+/stilC0oQY4qxEQVF
SWXYqJnkM+uaRoK2oQv9M56sYtdG691nIdfNEcmXIq6ZZBqqs3QqZCshPhvZfRGXzhmyjRguU1aS
ReWBHZek1S4DEEEk5oUbxTRnjvjWLwShkLx9CkFNBna2EK90zs9idqg5adVqe7eFdxoDRTn95v0T
z1qF7iEV4qCRRfTvxOBdCm+Ek8thwSig3idO6a3cuMMpCw3QHu7K0J+6OzPrJU91NY5On4RdWi6o
y0VmTuarzeDLwsWBdaKXVPcXLxV7k+CbJYtdXDWR5YvONEHYkKriSUfKYqSTOkkqca3fL/txgh34
IOx3kuGNtNIVkI0bGV324bUhaTcNcEB2HY/kDcNxAaAI0mghpFjaXyTFZBi3bOc8dR3bexVdi1if
ILF4uV3dUhowshC5VCJg92X/LC/2hskPtk0uzfd8xjJgHwS4kaKacn6GdebrCMP6V2sxjgZZuJ+y
lrvwRXwqSIb9i56DRrzWJZcJZjAlIGK6oWnmJ1xO9zF+Kqep6DKVIpjJRjxFx+mM2MF/o3LhFEWl
TSNAzesAyO1Ddp1vsyJDXouErHJComuM5DIB84UqKo4cWB+2cctdJT8D5Turw2wWjN2S1SMFCpp/
gbT3wJ82UDsBfZX3OFQa5H6SPzNYo7RXDzKhVhP8FMRqhOdJlDJ76oQ1YF6esPfoUYi8LagqhI/E
bvxilSF3EiEl0bqm9bJhstnSkXBgC74oFnpvtHkxcqm95b9gj9+vruFVBoz1SDtN3typcQOHD2Cy
PTQTgtLhw+VjP4jwenztBdw4SAvNpXFDU7ePRgOFeVQPbpUMUncAjWiEwX0QOfyr8YsAVnZtWZZq
gUOe7gxUlElp5odkffgafl5vHLm4prZF1v1C3DBwqzojRqbjyXbIizvnRQNvqfnksqWk2A4OpWNi
Uwmk4WwN+HRC3mLmgONRC8KhhtG38sdQabqw/nHueVBP4q1PncwFk8efREC2363zU/kPR2ilHc+a
OqLfsrFhWFfwQNg2vMIxCBlq5WZPfAhkUL75EkqITWfMtbCr/t8maohdAQhXYDZFn01opwlENymb
GUVK0tgFxuAQDqYWEO6cYOhsd4PTUN3+37hPc7kcTJ1UJCWf01fMFdRk4t5rqYy1npwIqVsoC9tX
B0Io/pTXVch6WkOaulSU3G5ebsWS56/nLlVTJkl1zvshtss1jZcnoaynuaoSVKhdSvIZE5q1JfIB
E9R/9TJZUxKDSSpY/MVa7+42aSS4eqJl+BA1CT55/B3gc0leg6dz5OCazYzvI3r4R1fRjgKYIGC3
br21nLE8F/zqzOIt+AxoSRuso8hq0PqnX8bG03neks62JDMsHmjO+Ys+rWaTcFUB84bq5iMdyGuV
geq2PeAWPcts9xhJV95IExBHkeHt/Vahj1De6GTCzziw++Ne9s+sPpe0RX4GVCoTTKrcQcO2tDkY
nDeI8exYZwvOaJLWkTRAxkVrhLyS0KA6v9q6DeRbQSRLFpY+hEDFUiSkw30ruTPz9tpfsjkIq2aa
J+c2YiFpk2W7iz4uJOgwaezHtjlD63FLwTOnmAucgicTE435dur1+ALWiuSltyxosyprYGsBauMJ
AEXP817fakjyAEbuhNF/tn/Ya5zHGjnOK0KvmDzEnJqiYu/DDPgPTLTO4P/W2eduwdpv9dEohsk6
ePYzR5JkhDW1EPn7SCTpOGF2uwfbLTfgdHj/yZEG/qo9ltOeCTOeXuUamwSXsmLIvUvAv6+kt0ep
2iP6xy5EIU4aTdvjwXarfLyKaU8WcPp1LKHyhVPt83yIrYjfjkVzi1Y4cPFMSEtVKca3ZAFnKttu
YIMVJJxcUSCtczLqWzI4Q0u9Rl7AVHJHT+k9cNyft1fZUdL+dNq6SPapp0E1dxqKKfP9Zr/V+GC1
fak/ltn4olIKdpcIE2kQCs8JCxIp9JMUfOPW5U4x90tycQxavIk5z4k/VptlZgnEVzroLtmc+y2+
cfpWxL0tNE9x77QbInLLTjgQb7bTKWJdg5fDuD8UhKnGs3PQEd5WTaiy6+UEyJXTHKqQxmn7ovAB
EAJiTQ5GrI0AwBsAu0xcGy+tN/OsF8bSVwkGwvqq6NHIbqi2sI/E3W3eKwGrkkhe7/zQKlanUs1O
u3kgcpNmAySGjJw/xHF8eFdlV/GfQxD7yP+W3RaggoJ2IMErmg8V5C5m5LplOIyYfatsfMk+TUPd
JwlvlpaktfIkQWbniMPHnh/IAR8YUz6TBMgZy4K7zi7zBKURsRUfdT6MIS4dpSPGUvQ5UeW57kNc
zkQdcecNaXesLS/ovMchpXYWX72jc8LsdMi7MO4L80SDmtLMThwfKoDRdIylNW5nCEzQ4x3duM6B
s998Dz0drKaMSPwhBWdTXCZjfy9xtdfx9BuRQ+yMZU+MTwG8+oVUxSv2k7F1ThgNfZNijZmUEKuQ
+q1CpfXyv9nq4MAxj/0zelE1tlXV/IX3EUB+/ttMP/uab71dY1HhCv89FRA+4NTMN+1nAp5sPEaV
L/X8vA757IrKIayS7UnrtW54/YHB02CwheVj4liMvVzVwpJCSiPF0OJo0p5HrW0siV0V2hm+tkCc
zSnsoKHnwSJDnqXLQDatZz3P6Zg/ySSmpvboC4kEzRliMMrdaKkuf99qpFhEB+7psdv3gqdiQzt7
76ph7XmyhP7lp96WVKsVVXw+l9LS1+1+ptuBofjabnA64btwIq3gyjLd3K8XDkltEmV8wQazbC+1
ZwaAZP8PhvNUyXeEPym/0n6ADT5ywvVqPJqG9rvdYMRAvoL3MSNR2FL92miUdiT+iVe5g7d2pPIE
zqe8Q5k7FIRTKnI/n7oPq/2YmlmhcSpGNVKomSxVR7bRSccmfd3REZx/UAKT8Oat0hlkAbYPj6ef
4LqKb7XwwRWhjS8byA0UXCJTdnHpyA7M3I/Tik58PQtX8IS77hPOUkLcuGTaiG1bW8Rz4wx60rv8
3BwGBNBPA/T+pYqSHSpc3O6pCfn6yGtszaL9Nri3iCmykkmmN+GVQ56BS1P9kZcW0sR2Y0Sy1brc
cARxFgTtxTJMxoQN4nUQjzVurZnTkhf3d7s0OxzrSb7mWKWDAgC3+wfIybYzajBgB1rXb8VUShRD
6gifU0+QMVozrpCtGWWLN90kvUq5AH6QRJpP9adUzxK+I8Hff5u3zR9LOFf478XU5+I3QwCRBM+2
89CmGoVc5EJkziYONQiQdQJFNmT5yd3IerQo4nVmYKA1aQGUlNrwXLA6JsjuEgYF538MvuTSR5g6
nUNz45O1DLmLk3BN4Cs5AQnvKvi9xvedHGA2TYb/nynseiF1cyvstkPppo/R+hW3MZhtZcA7kA70
m+dAJT333k+23kM0G0VAhvRs31KYXj9Q8t3xcEwNcCcZ6iQuD6rlAU2CPJJLZUvoPpnZq0sMpSPu
W+xQ+MOE9WG1IaT95rWM9o03IFnlY4Co1QtUeb57FGo6jS37jlkMCvXLJCxc7RtQcgmgTwzlADFz
8QPjC5D4SDxNVzZTq1dXJvJXIcT0W+41K+mJMZU27XNx2EjI8WW95Copk0B7UtvFkazLCuSGiTV4
Tab4ZV20rXvDPLrwnbYsvSovEX1mXjZC7uWm6wjPSIgT1i468DyzFX+gwP5NKncJLshqquehNXod
IqB+iaIRFKYE6pdRkiSVL/z1n9MtjaXgbeCGBrO7HcAlP6CXTOWpxKmmrEs45CLTwDFCNu9gwZk4
dA6FlaNs8PtjBmKu0LBSfG+VkdiwanNIIW57BG/JxyJwmbIHARIhYYe24ldvvMSAAhmMN1I+TOsQ
ZZBvAcMQ26if+/LNP/m4fxtBxbuJmZ+aZoF2T3rLPwK+3FP46SiwrZljQhvB4NsOfh1IbasPvY9M
pPyU5G7sNLamEz7cGofLrE6HA2LRp3kfUor5iiF79rNt+Pot9J9zD4jFIJ6LCauZxRwucuMd3Zi4
jhJXV2ri9D2jUeaB5wAovffRwx7TttnOalhfem2RNkuNLYQCRtjmyh30wauQFwBZ/3aM7F/cTeX6
Qjl9XXbF6RqQpn6dwog7odVolWjulJzP1gbt89ytZcBi/ViQr4K6AHwrDbZwUsiPvSnEAkjMvzrC
MAIFyevBErR6qQo2OGy3q5PV31AhvqhyFntnLMKQJeA41gwl2+fr4MkL2i5oKD2Cpu0Fkl4VY6jc
gPYvCr3NfF8NLRD75yEla+Eq1tk7FE84TE7VoYr6dvIh/ohvs9dbTv9hBtjzj+bT+YzpzUkSzZiy
4FHrtlmZ6sybFLpfWtWRecFuVzbVVjvWI4PPYle/f7GkIa6v/8XJmI9FfwHBuZhOQEK2Go2nmSAA
vSo5GWPzRWsPbuH5z4RdXm+HuNUy5hB+YW5+yfD6Yr3umFW6/VQwPdcOsuOeMGQfaPVcjoolU5Ha
H1f3ukP++irPkY/nwIyOMO9nHogtRc7aKrpysYj+TMjtDeK1M6NqGsCu7ybqKFXfqOInNh88iJGo
wblQ/McvHWHhl28mvnxNeBlSKjue0Nxn3vqkVgTjwd+kYDzGYfQga1vnWlZidtsfJu+J1rWB/wM5
EJ+ePFkKc6uibd7FYdbMuJbKlkNccryYhN/MyJYgqksRcExGEqr/KaZDncnSHTPdI19Jg6VbFkjo
sqxeRY4jcvAWANXfKJ8ImnSNTBLJFiq6NQk0q3b6+qx01RqoZv0m5aAqss1S0jMZ4YFyRUHeEvLD
cmqFWaAPYOLeHBUT07smPvKgErXFfqoAgSVvBtMWGOXOug7FJLG43KMLkEOQJ55TMrqYHQd76fRs
0RgE+ZNReZZPinvdmqNXopq2VnaNXblN86XljzFru7yemtcafjf7UQT7+qncHJkcjco4/4FeID6P
cz1Q0Ea3m18vd549vwHM6wnD6glwYAuQz8DMSeQeauAJv/CMTBULpDKK7SsKqTkLrCyPdxQ0qh4P
JEeVwB0giTl5aRLzPJW96Au0FVq4SvRaUGcru6kgLRdhM7bWeCAxp2VTpXwNPHuKmtM7NXzmxJ9e
hbVc4lJXcs/QHiIw80lohlo6YZMPesVzxtW6gIhruZ3+4kJKqWfhWwOC1Y+/Nob0Np2nc5nPtJW/
4OynxETdWeSB+RVBT9brTrWBCNIZvojICopZgIGAJs5ki9vZAvnYAfWZHO1QLXxdvTlS1FRCjxLT
ForDlUlXaQF3mlaCctbN/Sl4k1FoxxK5f9MoA90uE90HfhyItVeUSrMiNq1QoDyNqRpmIc3ESNeq
dV1O7AC2Dhv60MbKpNhHkI5FDlaPZBO/xh7Wi1lDlJuwTWMzm2tLywsm6dw04/58VvOMmPHlg5a7
9cjJq6gUMGGOZLmZrLqJ82yS0L6dK6+Q4ysSqOqPDyYAQ5seUYQp4q2qRWWBzDG7PTaJji0do1Zj
EtKt/FnagBGvbmuPNcd5V96KaKpvz+83T1oh6V59XGmOg7n6+ZXuNHrQ3T+gher4z2PNXOKcbLKV
+PBNZq5C48jO5zi449i1cSnqAUsi+BSP6PvTioNw91hMME3wA7MRKiwxXtX2aHp16LBZTzD4MrFq
jrzb/DHCC1v/L3UUzLpgTpYtfG+KX+u+uxs4cKSBL5cSOwUTpQbcsP1TEggBU111UFkKjEckK6B+
HvqRH6wJxYMsUVj7OTSy+3iE9r+rl290mYulshGVGgFjLPQBvL7r/nFhD0igTvZuuc+hy00Lrolj
7eQK9KVm5Wy1m2Nxp1NE6vzDKz12MucyihwRNYME9R959ubch4LyXYlcuCDvZxHoVU4bskJET+YM
1g0dGWjWo65GVAkrKiFVCNT6nXJqF72/jCsjm1T2dBpTUjn0IV3/Cid4O25pEHWwkLEYz8X85gnl
6V4o+qgsiNoz+E2AmgkbyZXWCMmIaFjLADLYiAMn9GHFfDmQ7ADceXWoA+JejlkWTt6bRBXBEQJN
6q6PcfNp1QIfrttEcqRk6xoi5eTouPvLoWuP0tUoJzFC9fk+ZVRMXUQd2RPMASiMJwG9nypz9qVW
fcqa6ZEXspQk7sFn431/TTNAAGgndrqHGdfppeyRv9IrgCuenTZ+JioaVMrRAikLTvep7JFzxas6
fsFbCFYX6i+2HVJKb5gMj/F2cGW5m4T6UuiKrnB0QLPxUcZTaAZdHuXKc1+taGVh4bSZ83DP4kc2
GXJIqq8MnQYAqHzk6UDn7CmiML6xjqD65bxjqZ/kCqDKB9iBpYDkLEbxIwleLULAi50e3DYXDZ1F
yzEe29aqeFHYcVV5k6Xyi9uCAliAqQGuXNkkq3gLRRXiGB6g1P9wWcWVBI/rfIgY9zAiYLUzv3T3
VNNOLs8A9s/FCybZp4km+q+J10U4nUSbsyF5/Q1ekMTIjg8/MtHfkdFXB+fEmWHjXAHBNqdd7lFk
6qXm+We7q5tS9BLivu8ytEMzHcupLP0AC6J0UcfN4axWUvBJi74sdGymtGGPw61Bi9HJ9L7PZqhy
8CrPJkHnsUqyhHNk0lXDX2BgIdbLQERcnaXQqjsAhCAxeOdxUpoMxgJ7HHGzxb8pVKwtAm8/efQS
sEK7Dy3lcMOXVkcdPl7d5deVXWb57pbqxF1GAbyVB+EGxQvykVf0CAzq4JI94c6cD6zoTmY/pVFe
wRw4kuFPkatxareb9rDV/01lR0+CrZsHHuw8vg1HGZtjX/M4DxhCDBVfb/oBzy5EJZ2Uufc7Qq0/
2yb+6C3JcgbLMzUTsp5CBKcHlxLeuUX2fx04n+vH+af5TomZKa773AHg+OnKlxRKkbb84HxAdKM7
wCLh7gt/QHhOFaNJTNLpRrcrSoOWy+njTFw3cNodtuCC+XRp+3Ez8MJpLEVMnBFczT2s09J/AFP7
CRZUHdi9JGO86MR8bp9tIz8R5okae20QmaEXB22H3DmDhrsTQ6RcXoEwDvYAGRbnEQEWXHABqyze
SxRY/3EsOIt4Mvud7NlvAoYdyF/b1jK2qEag4ZFcq+jwYmFTd7blXhAgY+cQO8Tcy5XkMtZMfKuH
GyV6T6jxhX8k+1jWVTTR1JXybSWUewZnQotoT/LFL++JBZgHhs/cE5WD0fuOiYo6yM7xnie2OSan
987B+Ns9sWqkG+TwT3Oht7VCNcQWxdKDK/DzxsMr2idatbJvdrioE4MWYNUWtDsihX9wNMhT/RZ3
P8/3p0JI2scVEJR/iTulIt4kdhUAHwBq17hgetphroZSISupsNIgRPczDd2tGVNYiYKMhcpOr4+2
RBUXhZl3WS/ZNE4SwD8MFk5c0HErtjdUY07SwNfUIGSqfi0yaeD9mNysitC9kLPF4KixyhHW12WW
y07G1/lDjD/sPkcYBRd0R/s17kEthH19552ExCCmFUxgdPygYnDGR8kAeYPt7jmerQJpT5IsprA1
ktvAtmx4WNuDt8g8trT2XDMu4DI+1qjLjLznLTHmL2yEBqbem0HgnDvyjOhTv/J6E0geDUcKJCTi
7lsO0ZQpaAko4jz/Ksh57Sb+XUJRyymWKGksrqqZFBj8AMSkxwFzdn/6cvWkhU3lzVQX2Wz9wAY3
x7kXp/YJmGZHJOeDypxxMfrT46rd0C8FAPggKm3Vv0A7JoGxjFmzosV2WKK2Bwy05j+ocmMpkoPP
Hn2/G2pFoY9y03K8WBZRwAC52L5phRqTFvSVd5d4dxbmRnXNR9RVTQIxKitejJwzqwJxlTXsraUY
6v88EjYAWb9WJbXBvpuCIy0EFqPnb3oPjAXElGURK6RuDBO2BoKtj03pQr9XVIttDVmTxfmRG5Q0
o5Vb37cq8iMYDA0r2Icd5oHPC0iWAbmB7iL6CzDVLsRTCjSTFRc1kaz8fgS+sg/Xzwges0gyasX+
IEctpSHzWcGR4mX20oOGCFkfovRhM84pyxZEuStkkLyRYKCrcIn4g1ZXRZG70xnDCahMGG11n1eE
EeG5+UEfjbyVI0euhIRvzJN9rsJygcXshj7M8p8SU0x2l2yFDq26QX8Z3GP/L0oZeT3m5n7neqrq
GJCyJo0fXdmarhQLOLFmCuAxfsZDUOnViOYYuf17YG60pDHVFB+ky0iKOUXOgeMGRoexVoFR8AK3
4EdexAOAGPZPCNsrEoSbjEXYx3c3uA0e8EzuYXwb2DFyfnKW8PIKmktdPBDWk6rCa0khr/ynDGMZ
VrPI2KtYck3l6loT5PqCZans0ul++JEiQ/tobOQGFhK2w0SVql4KP+wURdWfGjF0toE4rFZeToAI
eQdpVfa8NYg/LfvXYCUv1dtmIvweepqZwK3Vhgr8Zz0kyQ0Ed4Ceib4tJ6dwtGZIak9D+lTQ2bdk
QeeIBJYe8vY0T48tmcKhqWgTiHEz+wJogOc6cBC3diU041AwAN1qkwL34Sf/RwlP5zPLdvdzc7IB
3QwEDW0yfJFAGuEkgMGqi9v5lkV+Nw6O21c3BTZREz6EIhcOcrkbwWGpjmWLkyt8y7NXwCJuz1aL
6PIg5PWzk/AYkSj3VRu4IJAB1nsCUYQIx+bBqsf61id1kRK2pGeMK78oIyG/yGmJd+03H5jRfpxI
3IAtuGTE8B1/Wkdu7IpnQQjoQt18J5jska8o6O0jsyb4/xS4LRSqioTlDEuiLiJ6mNPfVlvS4K+F
3io9g0XtfWGmTRZujBUcbzfoy0GS5OeGVbsq3cCSS7NnluvTMXGLNdV/i9NrBpHiCOOYfegMYImD
2mUZs3ONFQLR3tD/bfxmlTeushTp03mhL4D1gHq5NOGMoJpVo6lttewzvPLwVlvZ1UKWkV8imyEZ
j1Cz0wa+Wlk3Y2cq+WCpI9wqMpn5qqMX9E6/kiSNym7dNNZUiV/L0coYspbxlwWnvAhVsHcvvtug
k+H9oTqNa8wW5fw/gWhmXD3gVqJFHmwHQmhLK7xVfJn22ifMnk7DnvkR7ZJKMSiJovlhgHM88iCt
SiIwVGA8EONwYjCMqKS2QFMs0XtuzZvWTB3h3yuSg7Hch6PSpce+CCzKJOlC0S8TXueF0V+x0zvh
+S6N8HHA127XmcYOxLtuRckWCecjfNRmublUFcOIeKpdvxeiOBOC1cRNa2fpGOYVsrCO+UulxnGK
fZFFmH4kPi7XYHG+vXsHcZlMkJZoF6XY1aQ0FRJPPkHy4Xfsi8A+mQZwkx49h2Rqqvtl3mOjFAlg
Hq7lFo5dVdvpKHWUGYkmmRd8vXA6OmLrDYN5MMxRwalLb1iuBHKB7R8MTzlLFBpawtJvzJDUUSmW
Aye5ATlwd2ohpZ2jfJ2vGGVi7/MSjsw6I5tBVj7ECKwhISpJH9rQnygCh5uZaXxUKhYVkMCFkVlw
bZ9fl0FeFE9dugntgoy5xgtG0XYsGNPAE3Kn9lv/Q6frS9S5yOYCehf97T6YtpwRwsbKst30zQyM
rCVTUE8t/1N6f0MwJA3XO9XHObJiQ/wPU8Yt08Nmu3XwOuJNs3ZatASUz222aspLSHSOJJEQhrrT
BadSqZw0SctR0yRRRqtplLeVPKHRx/ResKSAsBdtsq2K1FMJZJtH5gXOEywd3+WSc2pjBKdus53E
iyvqiUEmkKoZlrNwpk8etb8et5OZrRMGaHEyQmCUudpHCPQ4DhsOMmqJazZWOY8eQRjYSp3STWJE
eFOkMVBr7DPTCuZjJWDP8cMEWhpFQq1vSRB2joExmFdLQTtJFu+Y/RFdAi3tmDaCgNNyQGa+e6LW
pz2CHHFCIc9CXyAWAtAzVlVVjyBpJVqxGyS+wxccjpKc7ykmi7tY3fzka0FuNXwSvfCrGF5gmSN0
xt/qQZzDEM9CwC/NzD1IVC7b0BPPR0a9AHfbgHlwfhDyaLdcCow4We6x0+G+/pXZiZQXYNA+XriE
4xUb8fIeGbypG7ojy5+NjQvzhx7dojGq/70d+c5uZuKbXSHuMyZImIxGsWA405tCU8H0s+pDWBKJ
d9t8/7hXxJQdM8dXySc10gMUYp0dT8JZzy1Z4bMD5Il75nPN0OrHtlnAeSYfcbOLF/fG1gqJmQBl
I3/rkVvubLVpmGlDl9FahOuoWrldylFqacWoWDSGk/Yz0b+KsfZx1Kw9/J4l/r97vdFJdciMXXjC
N9FMdUAbOmLzBUI9/Dnboq0pThIw4W9hNWvwhFeJKVnXudvz1BBgsUyJgHltnbf+4HTdcvlj1fCy
fsaXa9YT6m6teOQGagQY8twLUUuuZbjRK4EPc/m/l7BqyszJgWpmBmU+zsMvTk5Jvv2S1RMrtu3e
pKUJygjy4JSxycpZHjtzJnDkBAQO+p1wFfQAKGGekXtV/7xDURn5tlJVmpTIsSfw34LbC9xo2RU6
5L1eYKq2rZC459vgBiBizOj8TPzSPqMXlYI4M2WVyh5csO2IVRvt7bJsbdXJFXAqcgm+nkSH8Hw1
1sGLiZnTNvFJUjNRHp1q/LA/dBVBFFxAW5wRMbeKVqRFbDPVYQyOT/dXf25puv3Z5E6fzu885k3a
uP8UEpewmHqkUM4J43OPGIDlcxuhU26IGBUb78d4O1DLUJHqV+WKhyvHa3ioCwfXwwfD+5oLach2
lE1qZkdp27iBqC9xhR95kdk+9C6EMzTGBGkLqCjlNcppoX+0JYaJk4VhJFzItFB2BsjFs/olCKsy
YVbmFwHMq3MWGoi/ptbMxnABps9dZll7tsenImk+cQhjgZV/AWqltQz1wll5cEmuaU3guYY23iRX
Oq4KNRCnXnNavz4FSbzucDGbni+QBmFy+ZcZhHKqfQp7S8GGOCSOxM8qAJli0wTJwkbCIhGM+a3A
v3yIId2ADAZ/ga7UP2ZvoW+oesal/DkPCOIebq7dLwkJygiaodWOt6Wd7ZPLP/tkFNwJ+lObn5HG
WZnGdeJw+He7mYogloPSbN/wKIDum+sbN30w6dL8D9ZkJWFERGLmhmfRx0Ndu5g0boaueoWi2w3c
IXpK6Kfry75MN+hFsVXMmqmUjwOG26HtD0/93Rwd9thwe6n/sJJMNmOkgxGWV512ldx6z65zmbRO
S1dPYv/dBvDeH96mQQxwi14jh6OLygd3PRb4hKejMhCvITxTWotKbZZWgv+uPNFPRgPVlXMXUWR9
1OSCFY8qVnTDE/oJTBRF17oK6F/welPZ87nwzCI+artT7aokNFLRfuJFQiNzGlGPYQozuUsHKQI2
dQjqhZ0+xDKuvizZmFGeSz1IuTlq4eazqL0JXKGsBbEPqNuJZ/9DuVAQlsPp7AjgbwD18nUIvotu
cUXpwVk5ap6P+weBW2EK5rk72a1cDCoAHOcZS7yChz/s/2eGr6Wt1YxJD/1tL1NIkQGu4j1uNTxX
Dq20cr+boqays/1VaOP2kA4r+DFlwUQTQtcpzjnGelT6cOIxrVewNc8PspuGfwUmXZkAeodcDaAn
TkUZQOApv2XkN7A2FCyoVGOor1X5zxixVhOzWInkyWsCheep6zfmQ8MQwCfRksvZWJNe5ICkiql0
C3hAuiv+tMem7b4vOa7WN9fjY6BlFnj9trQLiI6Y17lJpHba4xaYq0xHSW1fXwYh3LzSE9P5jumy
fs4WbId7s+ENhVKkov+zJ9FZ63/z11/6jFD8EmsTrjhsmNtRG2h4Ybli+QDGpJ9wH8dR8m7AIa9L
5pRREYZwjlaK9Xsi+oQ+Zw/GwUt4xnanoyedM5Aw1XVY41gtLaiJptN/lPiIn9hVk3IxEea6ROy9
HTDRk3c6v/nnkhbdzCJgQKGe2hSxFRHl8dPp45ZABimnvSHJTgehBDWKPt/oByP/6FzfvLDY5Yf/
/Zh7wsXou5EcbHsnhpiaHgKobBNHehbYpmEtyQ1ID0RZ7HXuorM/pGnj19ogx20az/zavIoEyEsB
H9VEgMsP4zENEjzgjogOzIUKNBSBOUaXNXHxWXrUBufWGoZxzUUWEItAOZjcgsG703NU4tc9xt3o
x6HyGGyPIVeze2/5t4Rd9nvY0SxIlnTucXF6HjBlCC4Jx7NPqHRRVmtEPTlZPdPTreiR/aNzipIU
Z0k69c+rAFtEQU69jE6QcIBr3x4JehMKd1jza/7izgYTYS39+rTSyRNR6iPsaDmHDE1rvQmIXGSs
Jv8bwsm2NF5/M0iPwdGbPoOYBBe+9rBg/w+SfJPvP+PcnYT3bkOZsA450Ti+WtteyVjnuwKn+bmo
2ErnVKaV+AZXtOgPWbVaBDpo8/KuwAw1p9NbrPMOo+JGJOL1W9j/shQ8OsjdM4vsNKBYdp17GXRI
CPSUbxsymzBwUKhGb3Fhhqr3PWSMleD7HKSCVy/ajmKPzKywnhvGY0/8Mo0PK/RK8ttFwlm9fDCS
/y/17Q7fPJlYI9ZwIUWZcB7NeB1PIe5vq0UdVqVhvSe/KlCPL+Z/LcWR9GRBGEUvOxIWvPvfvWKC
gNywj81iMzqdMnryqy83XYZ0lh24Byt+Xuw0w9/M+7w617OQbCzRWkWfEaIAV1KVAkkDVtjtTAQQ
98R2lmJs78Fo5ETIAUmDZwyjLWUfc7/11FWk7dE1TbQRW6voQzosz+9+pv0BRz8rXVpeNAsr46FI
nnbGUyMgLssz3gKwah0GZnQoeHG0PC/gk0sExnt+0IbBDGLIdRZPbVK2DIxwlrPVXKjaij4i2zcG
MPW4dlJY4RqHbDlSOhcDy1IHwMDiAxDfwpL0jhypEl0TPp4dBRQSnNhQHAOWLbyAxFeh4YIdG/kU
cnMvqXscLC52Ud0IfoEGRHZxlRCHyXeKds9pAhmf/0+h7bJK7va/5Jn/9D62DoyaYKlojRCxVjmG
G+upOe5GXKdmVbM9jY/JxCQZzgLkuhv25Uh2JOaA+37wSVxDh6g0TODqT2le3FneKV6ztSy4Tg28
bzteF9CqVLKczvcQkbWG8pKJKgBVwUkoOx0LI4gQy0gc2QA9E/DvXBhrhRfySsRk+L3uLa4ZYu1k
XEQ3lJ7tqF2ydsrV5p0wkdLEK6NDd/UD8Lh6WDiilpYIjgdrJw9qxSPEv5CjcgXV/LG2WdfXRkaL
hfV4EYhG1S80U+uQF4J6ArP1J3Iz5zww+2PTTclJJG0CD8X8U5mjq3zekhKPM2fpIFI4EzabtbUU
GZpjWeMfBGgeelkiAE6NXpTbpVv8nowyqF/VPWLuBc75Zh8z98qdBdUr/+ekx8CBtRiNIa375ZQA
Cq4phOElwf1DIzgQVM8Qrc22rfbU2HTgWAGCF6ma3Hjrofxu7AIICXH61WMtl65eUAe14q0+r77B
fS4OwkIUWdo/IXBJL7gyQxY/jg2pexeuiCK5DHcA2hxTHgd8PRQvwEmx+1YLuo6CPL4az6wO8e3B
GrqDcXz5F8HYIkea9SSR7qB3++DnlaJZ18lMy1ycmJe8oBNla6wS2GmQu3iapeTNnN/JUWdDH71N
jyiQTdX2hx9PC7Gft1waQhxe2JrWnLs4uq0WtpeFVw/FHNB8KyjjnEzSavLQTWS9pB+VNdn4jN4X
Uum97Blx6tq1562QMaZdJYpGjEXKAFQg+dKasavY7wHxUtTWEiAXxrcwUrudpHL34+vJUuWYw2ZF
tCKWJlr+SP8iAPga3Wt4YXxfMJrpQQpzF/VP9acaW4jgdShBQ3iK/Sf3A7+fJZMiTORz1dkd2KbC
vcMrcgTRtMlrL+8FwIHBlDfLPq1KrEvasBhdUbJ9qkFuBYUj/SPzmklfS5CWo5TqG6jei/02DvST
eL2T0To4RzFwl/t5k1zzKMMgsWT8j0KITUmYVtxvW9Kwl2zGt2OauqwgRCIS63srSGF+84yjp5a7
Imd2kQE5fpgoWElhP0X++K1g2Mss1VOrHHG3e6Byo1vwzjLR/tBRx0ATrjxT80pvs52IxUt8ueQb
aI8F6wdZ0ZWcUuwNbUCbNzmRKH1SQzDwNlT3uLiAiyohO1tWvPm4cgQf3Agq08M6rihB+qXrf0zz
w3aI/CC37SEiZ5Z28XuO+LA/uuJrpdjFJNcgAu0OG8jbCL2rr2VmLRrFB8PTconfrYVJd/9ukhxW
P3iEEVLw0ccDVjoEr1zXaI/MvBoRCP15dXaWgkXOKapuqxkA9lHJ4bAo8YiLGgLsH8WvZ8KEwhJP
DNHT0MqCHKfnoKUZOjjoXhcHLDmSTR+myjQLF6cDUpekxp9yXcJSeHW/2kzyjv2Mw5YkLOQLv9cz
M0FW5QXtR2Nwyp2QvUEO4tSe6++oVteCOf13OesdadsUUdIfqJwIvfn1jLT/4UmTzzvnukvIiyRL
AZNi10ku4G4bV42wcZPiugQigS2vtuXObEZYkeA8QH4xzgAMFNjzYtKdZOBHZRAPpyb6CGSBBmda
Fol9AexL5I5XmNBuKI4WtJ62JtHJKkTpMjAzgn6AieuuG1JUtbJjQqJP7XVkHTSQOnVNsCnfTuTO
5huGGasjmekuNS46woVYPCii9RKDv3oBcrmA3/DAt49ynx4jDPQKDViGcDy3Yrb/T4wf8+ddtwCG
ebBLQ8iWw8j9S+E24FGuM7jZ99Wo5ZHJyUDZndx/7fMMjH4G5dXLbMbt1loL0usFarH0rGV/O8U/
UqMSt/i+s5CIuC5rEVuOPudbIya2w7vRim2bBb/dWwWy2EK0NblckQRbP9Vg5VzLpIrPpfJjeN8Y
G6WEacCB+fFoAanapuzUkIhhlu0s8rUK4H+UjaRJHpKPSF0ayJRaFhRRFKk4ZlcoyCltj8rAcmcC
bLg2bOZw6OqvQn/sUOfDcV6AqomqfDgKMSmv3IQACHOZZqp/9TwqEStl07F7QbcEl+1AZSVVLS5Y
Pnl7NObEMK+QtvpqbN0klhNxVNdfG3GrTucsBVEDbnIusaiLXNQ+F7sNd4LUwboKGFxi2N8yjzO0
0FIKB8RDpPx6uATxyzaXsk7GU9+jlMV1tyBJo9mwBWqT3oQlNpMkqKBuS59HbhjxSwOzrO6rH8LU
PsaUPhaklOH3CmcqickmMvIBwMlk/h+sEk08jiRFdz+xP9NeJJ4fLcVDF9h9I7/C3KajEK+dIRs6
6jRtwXic0Cc1p9Qv6VyL4vayxZ2Uu3UtQE8bPB9TuNS6Jc54OAiRRwZZ4VXgleswkbR2kpgAvrga
IM0OjCCJTWbqPJ7cGXrKmldW17+523eoi0906saHeYe9DvABx399+xryxJ35q0/45KhK0ea+757r
3kOqze0eu7lAET0uFKAWbYf0fw7lR8ZOM2EID1x1xXc1ZOE2pIK535sepoFoebBiEpCc4F/WSjx0
mO/jEfSppH6VLn1wh1gt1uz52J0kwMj5DhLV1v/FCXX+DVGs4qA1x2jznu2i+PqUaWKmSo0lxolE
9UHKt6dkJrvvkpMiyZoKWF4YqC0VXvI2P8ZMnt0xfWyXQNCNF/KovgI0ZxJj0AyfZngq/1mpNeJW
OCEAIbFEyqEvgTiqYAvq3YBhKMwy9kirp5q/2kAo9ImSLIz0eeyfASjyrQcil5TKAYHiQCn2X3om
QWzuHRKgr2Qi6bEXBfjn5okaA3Bu8z+31bxRDMcayV5m2ToWuI3Snwjc7XNz2Ee1ycAJz2qZQukp
Wioh91PDHVHam31MfwelMOVHW0E65SlYQ89SK4dcFYchFkCJH1CVQcpRf/UbuVS54w+W4UoFlRTB
rLgzM43T+19HOj7Dff2vj66qG/i4nZo5IH/GeItqOpiu8+4mx4v8HmsST6MQaoW5WbxC1o01VpU+
Ei/b9yzK/DIF3Mt9H6564UL44c4TYrESVrrQ5JmqHBvVvEp/cbCD1EVmfTAStpgnlayjJkuPQafu
iByR3FDMON6AY0uwOc2J8fXSN0wtZXktCJ8Y2X9o6I9T8RwqEL2/ffDQAih10gn78D3Rnww2MB5r
MfoObh84nfpHBW3QjLco7KlkAYkCBNpFiPbaWvDLQKFLCptZsJweBgMacZoJdJrvENcRSGRiIC4J
fAAMN1hgliz2XKhxL0d+I+fECpe0xx/brUj72Eed/rrMcSC3DbYat3RHUbWEll34ppwm4BGfMuAA
TarZNeX9rJVTRBZ42QFytiw95Vt9txgfJSlMMaK5VgRMdpgXr50Xkm8ZjcGdiMDFGGGdNrWSXXJR
mk0NPG4DEd0VLcACWJdLlACRnWUbxVkXuGfxphiYJrPqZceKXNAHV4TUBH93UZqh28mICubF1mm3
J5nSq67+e3Q7w58v6MTVjztJBCzNPG/vA3P7zuyo8lhflXNK6RVMgabjhUIKKokUVvUXaoeE1JIF
iKDLrVkhbP4hxxa+bUxJd3C4LizDTO1mR85kmWH/MX2RIAGBk+KabHV2I1duaPPr27hhmt1GE7XK
0jEdVLKu+N+rDqRJx8DjfW1rS39fHNTNl0UZMmqvksZlszKftniSMQWq8gSqfmReE/a0xEuZzgNn
oLxyTEfUlcM1DnHeblrtaALoLJZAKUgugG4evZ/BaboboWlZ/N+x7jAhBj/2Dcb0tx6CI9Jk5bIE
KGH+6EdPghjZgQM+0HJDAkZJ1HeaEdJ/erv7T/6U2s92akYYnGhhNrQzMtw7EzbD6bPTFZM2Ukcn
eqD3RqJuTBcWzb/+qbrvLTs45gKyL2XnHcsXCPTztwGDZkGshXHb69sAK3Hj3K9e0fHN3CnoBPf6
IzfmG3uO9K/6s5E2SbCmO6E/PFBkNVyn2bncUfsiy6FydJ/UGxaYjwNJTTSHvVv6zmU/H32oHeOw
VWnVC0bjj026KNLvwmuAUOA46r0romJjaaPPSIQHxdH8Z04aNqS0uZUVrHnky3r+nlJA9m2FwA5i
ImNO+V7m0a4frFlLsnAqFy+B9thrBLjjc9+n1xjW5De59ztHs5ibs47OcZRqzMVb0dRSiVVsQBGE
/0aVSUPfOAB5sHsok2OIRPCQTRqedMqblOI/DjwgJMsKdaC/O1NIqAeNkEAweCdgc/03VR99LKTm
wh215Px2TrujlApfV6rTOxNAYxlXQUxK52UF3xNHXjqDttAfidivADOZi2Z/mIL3Gkdk2eUxh1nE
I8d0aMvTPZDwQZcltfw9JXM7+LVXSlX70ssUWHXZOi18Ok5dCN5sfz9FMA48uf1vdVArfqYeJU8y
mmkfVwpj31ABIJSiynCm5aoVHGzbxfAhNMu19BV5iLQoJnkI0ra9N/JUwYfJyfvqyTdPQhG7DQRS
qxcNzbK55ThNGUT6HFazruVSbdAywrbS1Awx51Z4Yuro8Z6B8n+/GInLL+UgqS/cwoN3Ed6WdCL9
anBxrfvzh2n9Igqqd/NGxiRFQq4XDP25QduT+2ymcxIHodHMIyaVPrzSz2Zn1qwCNTDA2gDGW5nr
6DYws+aOOMfFnjS3/zm/j8GSiG8F9nwIaExE/NSv4ijGEX75M2Ao4zvgSnI2S3SJyeO9oxswX6jF
8OKqVNULWk27KRp0F5KjlJngyaeg+AogFxfp9UVoZu6OGHBcn7V8rUPhnba2ieXrEtA5VkpTcVXG
cCffl1GR1U1codbLnUv3uqr8oU4hXUoVSwmgXUvQ7AGOg9fv9W9VfYODJ9xBibyxwBb8X8bJggWR
MxFP61Wawn/2/FoK0fiO0BNA+etZA4P40PhRg2wEyIgc6TcV6+FtHBrCwtWreD6ZlqpV9IcgUbsU
OO8FIifbd29kmrTfrlOEX0PJYX2v8c0OacnPqjbWKY/Y9SCmhRhPkym17iNTmUOn/Iy+QBJ/a1+m
1uoL2EsdFyps+lF2cIw6HjUa7Wb25CTdXYeyAA9ODq5GgMlSBCnyjuAjt2VslkPsHKn0FWbzlmQL
OXRbQTjbgsmYoMbqXZu6x57FIcdKu1WIeVT2XQsdwgXTQCpFFFnJru4cwQKB4u4o/hHyzyZ1jRVE
FKo8X0YJoka9e1fTkYpwasVEIDXREYi2fEtEg/jvQuiaBDDmrYhGRxljnxV0NpRc8NvkxqHwQ3c5
Ess/3CEDIrIaoGSn7gcv9MJcLcAviUVGx33jTWRvd1Vm9eGycJMs/+4IHlKVkWAvc+vjyrGhB1jN
NFNTzpvA9N0V3ITVNoL3h7ZOL58OXSmfqOTaWHRXsf2BDggyhqqY0S9H/WaG+19o9L1cCXvU+ceR
qq7tV7ctiqbCK9z16VnprbClu//KvMRFLAta360p+G0vOm2TXU7geT0J+PaWW8u/PYs80yOpFuzf
NaLLaNg5odsiH6hM5YSG9T7NdEswwryhFo/Etd5omKcUQxaMls7cAHT4+28L0W1huUBgrAXXnjkO
UAhg/v3D1xCBggv66qcAmn5GzJKxHOLkttaZZMDTkl3ch4uMd0s77tILbQDr3XWf7UMwwT5Wk5y3
dZkiSK+hB6gvFQo1NUHohJAPGOiifEKIOutb6WKK0s8H31TGyE/vwtT4XoVer4J4D98bStQvYiE2
+lv9N6cEvdIfHInvyWH7yuGrkHNvd4pTPEuhmTsIkWWp0Hd/PXiBUQCVQr5gnzT/PocqeXAaHA+o
/tgOlZXq0l1ZyG+PCU1dINuGCh7ywd6TO8kJp4ORRuM9+oEEGWQ0TRUf7GFV7iRgjy6JlJ65q9jb
XTcVnFtTPp8z8K1+0k77gK2jI3JxB6sbAg07SjXbT1NeOpPGFbmSXkb2ATzw1ssFPXKsvuUb0bKx
raaf/mQFsRg7txDo1rH5TJg6KJUtMcBS6r6abJmnIceS5yYTek0rNVjfWD9vKVcv7W2wLTiC8CSD
msKtvfcTQ4cCTL6x403uX4+tYOAG94ScTNpqom+IW9hMKy9m3wom5tCjk4x3B16mmrKNjQulbZQC
VBg4zFOSDdDweyQ2SZG9HU3afeKZNXy4m+AFL6OSTX+dSp2nGQgy0WjnDTWzqoqMK9k2ZL5H2YWK
RM+vJ1TDp8suQjPRdqkpYnF6/SfdC04eK+FO/VYaTZGC0sT07n7iQc717IjYHLdhVfO2VMZ+WFBA
81QYx7SCZWQTohScblmyoLNglCR4qZWyGHgRCcGOecnQECPEWQV1OK8eJICKV3sr4rD/iBmpj8T1
gK5Z4O8zptio+5IDkG7AI4f6XR5mjGSV/Msehpi2sMPAFx7L1O24h8L07jOMDgmfgFffFcsfDSVA
W10fyrsbcaNfS+TTxqewpZEwY8oh/mjDM5LRf8GUPVLs0GJJZ39YWG33F1f2gQ6n10tvgJbSdmj5
D0iqeKeVIgQ9JkWLsrXHsl2x3Eoe3kgTvxzVJub6t5oTjdaPQ9ksK2dOPGw4EqdppDG6nHtHvxhv
p27Rky/nJLXx2AXeFff2sRpsjycutYXad2249EMA8msPfqBMonC8hkfEQ4dpEaA6UhLfvHfHF9nV
tDYYcHT3EsoOmyNbkUgKLPG0ZPI2aR4O6yYC/lQERpqfALGG+NPfWlsCITUwZOLZu2tVZkYfjoEk
HJG47mWhAzb7eEsbFmt8l3Lvk7X2itA5P6Ce3hesBDPK3+KaIZZBA6/jY9B+7MhBJFDo8cP4XHsl
ElrmZfDTOKD7wSgF278kFdNYh3bVO5Xpb8O3yhmzNsbQaU8gi+zXTD2+ESFYdtdW0NIgV1W4Zx6W
kp/BtulUT20hYnsdFRcrLet5xcku0XoZi619D2eqvcGRqPyY2PEbtKMXiRycaGnNngFh/IQrzI1j
a0qDsHYfyiRbgwAIRRlkv6SSPi3skL/X17CTE1j+brW/HPEdeYGz6289hrys4Gg53QFXATE45N24
9BIMdKq+BRZhPNQqNllgQQFxQf+NwvAvIzl8Kfq9w7xeCfOYxUd6GROY84PNFfwKlpvAZwBlUy/P
4UeCCTM5tAHZeHqgPkYuJaN3/tIH9YG8+tzMAvJZBKRSvOJsKE42uR7eawb0z8gZpvX3IMj1oWL+
iC+EF/UH/tnsVuWVWZgMBPQ8VqBqpcCLLKYw5gOGesVzAn+Ybaee8EJjHm6DUvQe0Wk8d1Gp1Uy7
Su1oXHG8N+DAzafL+EqZCqnBsFIs2c/XBBWD7xCrDhETYEQBdHVWy9XXArPMxIV9Nd0HVEsMCV7+
RRQH6howPfAjXfhXzZnJPTDDGL5TrmHhhPjiB7v9zicFPcxHaOT1hP0lkVhghXKLVihEba6ru10l
nq2/uvlcFsdqjatJRBY3ZavwQKCb5iXQhtS4U3MKRuF0uPlsuZ+TD4Skv9fkpPZmngWeAnijzaUF
9mFHrqiHis2haENXXWidphNJCQ/loIlEOV9GdjHmw2g3Q0OtGD/7Reb4oHbwYtiPTYc5hwo7s3U3
v4/zaZLFYhvBSjEPVSQ+ic8gWqyk09OVFObFVZSQLDvdNCn+s9tOvNEH4Ba/nm0HeEMLpbLti41N
QqPjRTPx3rDTBdYAI6R5coJkJLGIRJm5sn5qY+xfzsMFDAVTz7GHiK+faanK/2hg/X7OH7uRssJ3
Bdp3tqpaX109I1S/xxXG+0MrRO9etGh+5LO1KrE+XgJPXtzYVffZnbO94c71g7h+4YsOvaBIFjw8
vHKFW1P9PceBRIrgVuIfASWAejnRZ0BGElmN9J2DjH5XbscqfrM6wWfI1kNSfr9HMm69tVHlQPM3
zqS+rUwkNGgd6S8ZVeGp9gVaY4d7yVm0G2xcNxT77aCqVVY6NWKZ1dtfK09PPp3NR8F5Sjiqj40h
I7gMpS7sGcA2cO6L6DZelUb/MXHuMJAqeJCZlVmRQUQIMoBJBM6l7B8dSYGawh8q4nvYljJn475X
VvXH5Uar7UVfBVR9zHB00AaHEqLwQQAsZLdngLGLeaJEC++5D3AsnxL50jUcyos2V7msoneA2Cwg
USXpGkI5EXuEx3shrya+s93qdimy9P3WMVWnhr/Jv4cTM9x1fPZyrQTmiRcLh8LMhwW6WSAkHEZY
dEvcJouGE6VyXvjnfEaZFXxj8dmvTAKz/0AJkAMPW69+ibr2mZOcQDvJlgZEHx41lPCQDfHqFkor
Vmp2xJfS4eXnoAqZpP9E8ScZV2Corm34bP5ILPwQAxZ6tQs8uNEYnN+kWIFamp/NOUFxzLC/FHQi
rn1yHvvLpWCIP/wSYeVdCh0pgMlryN/betpv/MdAtkGkZ4nHaI0V2VBMYdiZk6lMuGQKh+nixgMV
oxeR3EMcYEQeaIv20XB4zyunf94ztq1QGceSUBOKXDpLA8nweBCijrYMBJQk7dwFho8ONpfudbFD
/FfdqV2YXyhWvxx1MarMbWLtTcGOND0gysfFmM/K9LEwrQ0VGTY83SK6qoeuH6dWuPPxW3bqH62S
LllCIkAaBlqyzVMbWP/DT7ZmNnBo5fTy1cVpqP+uAfbo0F/HwtqLeZ+/svgJgEo+p0KR2PQqGLsD
r2BwEAQqqq9PPj1J1RW8pAZZtjr/r8ilmupIapUUuztRQpX4eGwR5jhBQQJ3OnGy1S7eQa594KYe
PCE+HnXODI8Iv6h+ys3l+99wqPv9y6Tjw1OOvwdUEpr5a3vF5sCyYTuP3cToC/Z+N3K/9SkkQKuq
6r8Yt5b0jIgRkzTFjZHPj/cZRUI3cmXTgsLEZNdwe+HbS0QsTnGJXUarhv9v2IIfX6Pbf6hSwfWz
VAbXcXexd/PFu88CoPruFBl4eSJcbI8gSA3GJzk0qwYIJo4GNDj47Ex2oErQlN5i9KMOWpzrGr5p
33Of4L8zY2ogHTTlLOOBTEe08m7f5hsBi23R6yDhamrdqFqjoHWppCzPJfpROVPcWF+eKAAg/9OM
hbNxRP2F3sBa6YkDEu/T6srSCGwNnOhvA/M1+HV1ywZil2qoC5AZlmB1/Q6o9JHkUZHBwcC1SXCD
TldINHtXSXqTZea63Ilf1btCM5tNoAlA+CS83qzZ9xirqU8WZO8EvFzKT8e90qRaIa0aIkiKU3R2
1SiAYE6HOf7MY5kgNcsKkLjwJuXisWOKOl3G6ru4MdhobuWzf3HYjV+8CuY1ehBH/uEfFiZQvkg2
H66P1/4kFZUciiBgChF+blU8HXf/WavGo4xRpoI3qsqAqTXqUsKtIt8gEnKqredLX5uh5dyWpxNs
SKubUc0rgsDMwnVOjHCg+7ecggcmKfUkbe/MDGeChvA4WGy3BSkVDw0afkhZaX1YdJTwxXa6CUG7
ktcBvzCmGDOSw7yj+aFjfvlP5WQ+DR9URDRgBIIMLBW/QIGtvU//zGwt+rT8p4cAwhJL3g3vCUFZ
xJSDxpp3yZv7RV4LMn0JYZWFF1l/ncqygkxklbROSWhk8v0h+xo9F2NH2eyiUCN51i5o0dt2OYeV
XsAIFgI0h/vSPaN6FOA2qk7noxz8WkJ5upgcU00FX3SoBk1f9PAE6cKq0kQvHN4HRIgVzoS6hRks
TlXBKKkCSK7T58dWVHAmDokQhKWhM3vb5U4MOfRXa7qVEX953UUk6JbSKbxNWpH2l6tb6pVNh+ZB
4lM22kjhLlsriY8oCE9Xrd2HMh53jmbMHaqbAIi4mY1qvcTm0Vf7kRshZzJ4VKCxCCxQ8pl6B8uU
6eH0g73DCZ7BkWnTqQGYDHzODQuKc7cA4IsCTf3w9tXbq9w9oZM+8QN4aMinuATknr/ZAjJsVU/8
EFLODQdQzZvE/z1LBZTOjSJmNc11PnF8FLuqhDQM67j5f1eGwMsPa9Ce153oKSdtlMBE+ckeghWF
1yjmz9b/zFKS6ZtT1R10FgKRWzu4xwEuTO8yfYIoJctiOixt5/l4ugtzt4Z2xixbTbasGSapc5mc
BNDWHxlSqnxmpUg9PS9Xh9LjgVgxC8nLORGHq971nevgBg2BNoTb6g5LI7X4lOfFG2G4glrWlt6V
74MzRMWIs8PqcKf/UDL+KwLjfAstLaVrsEKiY+ODOEG7KhIzNRTWHwbVxmDl9sEyCGY5SicfdYui
P/GwAZCUgWtkHKzYBi1F8Pvvnxb5z4ZeU9gUcQTaKI8jvW/IWlNY6gIA1IVuWDDfSPrRAZXpIM3f
ta53t83tcglvsXq1nGpOeL4pwwMU/JIBeefm4M/sd1aBj8cUjHaGGQT16TDB3lLcsTRYfTRBqE4F
Ol+CISTa3QeDS5Bnva9WVeOEPJe9fCVMUVcnhz733pyiCc85vZalgjF/v9lBe9XNxTmhHF+VJh9L
TjOdMTS5aNSjJ0lm4Z2exPLgIeWrQwBtpLl68V9QsM2zIbKVILtqUbFiDJHNnTId0PHXnF6wchkk
zDCTTfUxtsIkNyDJ2i8ui99OQ/eUAl61TGzQGTpqecynXvsiO+kjRg7+WAagsqVAeR4Mfj7KOTjj
2CTAEi9oLyJAUAxtIULbGgzNoSMBmIKmLb0C/0dCczgk7z5mPZXiQ3e2C4ykWA4QHcaC2qJ6izDF
3D2QqCkyqDDntPjHwjxkqobX2xaV5pQ/9bwxBUglEn95DQAQvV1dmkhjQH2OnJRFikSMoxtaJDeD
AmqAyUCCOBA2aXGOtvLeSmvVQq0bWcyRTcTjdHobehz9Oi3Cku73E1kNE9HSSSSTjC6sp5ZzFeir
SR82I8li7jdzEr836s5xY1FfFUMRDu8jdP5Z1UOW/0IZCglPsiC5ruGEyK1DXDiHVDBlLyadGYfh
g4sG+i0R3wPpA5JnNeKWr8wXQZzR8yed8XWvQrf0ONB9pbgPUzI5YlyQ8OBjdMct3nFdJOpwETan
ZHztkV9iGumJFgLZl2pFSh67rZjsKuuLt5B/k0uinbvaV0HE6MpXIEqOZM0Y4txIw7XEN3bv2mdZ
bswgDYCiBkL43Ev5kDnaYmyPNFIVvTpBvEwgoHCo5F988BcSx6fEYPQlwtZURiShPb8ilZpJL01E
d6hmGFAEtJyLYgyE7JHW6uPXQq68JAMSvTajF4+FXFMAhrwFPaYWBcPR1eIJthXZ0kKGBaRyYabY
qfYoo6P0af7EvvmOpqKmX0sj/N274Wm9jt1lUWg00HaJVMZWJtcIVGHlIsUXuAbSghoY9d9S89ep
DSaV7CuxWUi7UYANEsDVzT+cHw+IWztm02Q9YWDBcWvsM0/w1nDgg8Ml8mzFJeZ8PkSVHxJChGsH
wCFPMBF/kwsUGsoQq7iIR2XDMX7ywnJRrfEPOLxrB00lh17d4V2Km8zguKZdvGyn2anXQw8Z7EQa
mMdz2tUiZgyCQMMN37QrOQDeHAHMpB2Vse8QFOKlTcnP4U9YS7z5KSUvv4dqKX9PS7Lj9yDvMAHT
ZGaCWgQNuqDyO0U1H6E+/iBQBWrjf1HgRzhMXNErLqyd2FlfCR0T3FjMzl2DYkQLePrgOAlWY2s6
qrDCuSuMQDxRlQX1Vkgru+izus/EgYe3f3O4k4rFYrhnaUl/jb1zmzae+CY11wyspYNgh3gf5Ni5
YXVALiRWR55ivw3pCK/qsAq4gil8JH3o0p+lQStiUqTEnEvWz72k7RaUJr2gPmec6j5FYPijB2Fa
gfN1vsbME1ZmigW7iMbXuCNCPoNIQ5qx6HrzyeR4v6sfIihXz+HESnITQR67wgSdZYFS7Sg6ctY/
5nqAyXZcqVtl2gLqmPe1cxwq2ZX57EY/MtBpsXHq45ouQ59JSKbwtfBK28OltQvanPkZNztZl4d/
qsk5LMAiw8tDqt5A4XIADNhSJPrauCXmCKCeOAvVAP/Eb8viOvii3CVfY9HtHsWaQ9efya326pzW
BbLZJ3+OBLJffB4cti+Xq5ozVUITva3qbS2vLc9f7iIWJoHoBQ1HRPrRr6GfG4SbKNht2MN0jLnE
Q6w8J9j1uxGRkLtvfzgnkvXMYH7KsEjzA+osHSYvb91RLcTDOA0CLawW+z3YWwQmpRmrQRsqqWjQ
K4vmn6N6kZi7p4RXuMnFgJoLPKRvkbyWbXO9NVoEFT/gy0RtPSY+TaOjK4aNgWT7jT/aoZhjpIHU
qtusq/J0snax5l6Td9iU+LlCN9HdF2S09z55o7m2Z78ig9ze6YDpmXuYjZSLTCMu+I46/6sAy1at
W3/Nja0iWeo3j+RvER8eXv2eXBfelzvDQIUReZuQyRBwQ9YMDwXoM6w2hsC7wmeEMQIPCs6YzjmM
d87YmwUW0vNw5uehMz8vtNF46d3viLGSLpMfrv1whsSKBs1bIdrqLnx5rEsNnHXjZz2JuyNVzP6Q
7pWdaf4+P+mBMJduDnPaDiULMSydWAcY6oG6kPAjNxdNb9KMy5vloXghbUUBeTib72jA9b3ZTDeg
/a9yhX40IfG8RbjnsMMGPhrPx9pwwlY9cDD6xAvoDgMxS5NoAsA0iPrTwg0ipl9bf4h9tPyxaB8P
cn6L/i2oqhc9ZprYl90QO9O5dmiOj0cKETbSs4HaWY8PbYHUwr4vUo8tbMO5Q/a7wKxl1TPWhDWz
nb0UzfM2oYajCCzSfzlwlnxABYVL7SCKOxMmVJRWG90O4Imt/hag/iKvFq0W7xm5RSvI18vdKtFd
N/xtNRuZgPl81Zosfjg/jGem/tSkpg28K5nwV47fnX0knerKa9mrUYpomsrZld0Xm9ovZ2gQR0yC
FVhCyvcd6w/xDr0+sg0XpVNpZyLuMZSfhLhZD7GOnFQuSbskNIW8ue61fg1HtRduiHe3Rf92UtH2
9WUgJmYl+CCVLQtBfV3OLlzxq/EC4lqwNYG/k8k23JfGCtzMOMDNosH60jHvwnHnVCZeU+jo2Etx
kh7iAIQeZyArYwqnLv4Ialq/m4BBqZlKmvPhnBOQKuhWWbdl82yldTTRwhiTKoMnZQS1mT5oQw0Z
kK0qUmX4iA6DvQYm+ZeZEfkY8w2lpVwBlLKAn+Mp96nU5xveZ9OTM2wJU7T/F+3SR2tdTOF4TYsW
qAyKxN9kL5xyUavZr+faJPGwCS5QydsVpmJbhPDG3n/2Dz72P6ngB8Z+/mveotDyxin6KhIepeLT
OyFxi7cDkEFeWYbepPdetAUcA4nuN15srlF9Fxni902cnCh4g9nASJX9dwb1Jebfo6vvxE+LL+l3
ie+MrAYDEIrTWJ583yTRZH/elkUzqd36IH97JcbzLiUHZyv+hrNHU9JESbijFrmzlAX5/W1hd5lR
u02woh2GW1L4eb4rqGtZq/BiqLJ7e5+X+HzCb2gfyWmcId6N7jcdyGqbtj7gnOeq4810mN+5pMsC
1Ucm4kcU0c9teHW4EDbXCDhY/lNtz5DauarZZAcaIj7sEjz2KxkjcTSqlv/8UQKuwDervolKxru5
7HXo9Qvk39rjcCZpSI63gZ7ljsLWeteOObh6nBruXPuRefUEO87RwaWXxbus2Rg2DpUTRB8vncHg
7vXVXd9z7UmgOC1LdIRdH1mNbokZ/wPOTA0yRCGrjwddV9TmnSkCy0I7l2QC31+Zv9jt0rLAGKC4
ZQKbLkVxQGCLgpo6NejcZUlbnFEmOlB7JRRvmkjB46RtwB7J6LZi+j6uPlbL0uMxRT/7sYKnnTcy
5xXb2Q3P3FN8QMGOcGIzWhnEVqVUsJhvkJh1LcdXmu8nkfAS/f4mBZQAC0duKSKiTzhioPzFTKoa
7oHRjgqQWgEqAr/O7poF2vCzxzcY8eSJowcqYukoMLGKa+ZKS0wUKuhubCtIa0JTCEs4gzIpLYR4
AzCeMUWbsl/2mzfgd4Mfa892wzOBxwYik3bWxrg0APdy8IoVV7zxKTDUVJ4I4V5EufVvQJNSGLNW
ivx1cIOf/RtryXVvXnVtTJjnyEU0p/3Sui8XInOXUebNlL9Tw1F4oHcOzTBsy7IUHkBxcUwthddE
o9/PC68txasU1O1YXJCkXEef0pbfEGPjSetEEpUXi2MSf/1sbc7gNg/XHwhgH0X0Ii600HPq3OP1
tJbqabEDcVBVi/KcII5EJQIjj0/lcFcNvMLiKmxP5JL0Rc3glpT3bkcijnoSRII3l5mwt4hB2aD2
fCdo7JfuCK0+SDErBqgg7zk/bwnQ8VTFWMKSeJOnWmEWVqnB8xTvnhCjPTc4t5CJI4weTnjjvGJP
GAELaDZz26pJR3Qn9EBPmORVrF9xZG6s3bFJQZ+zKY7Hz8YJKlqZaTz7f7XyEHQgLmrXFoay+n+G
S1nD0abZ9yRbJBgi65amsnuafpKTnFuOYls7TrW8QuLUafPo7CcV3zvHg3u1b0o6YV0i+4w9oSRC
A1UbERrs2szNrQiAhZPISKHZoWJGY6SdY7SxyYAl14tYLSvCHho5PpJeWbHmovjFqAo/HRawnWNV
QJEUG/+sgYtvtYE3YIaqePPjnE4lSkffmfvAOATuyK8Bby4JcYT42JidzyRtl4aEcAnS1VPysmj8
q/3gc8XfsMAHCVDtoQmK2Sn3NDar3R1PUx4o6QEyP+Nl9ztuYNJqSSmT08EcO9qMMICIaJotUkdB
F8Tnb4kriCeEEY8JtZfP8xe+IrYenfsTmnA5equLMdKrHMrklM0RfdfkhLv6dc9VXI3nbwGBtL4I
k8UdeXuvVVFAUFIS0O2A6iyNaSnlO9qsVGGuL9NKx0fVXunINWIegDZPQClYhUXonzXrtysrT1hu
/raGGU7JSp1m7cfIsEDReDtqJo1RdrG0LKo6w+J5nuFI7nm6kKf8bVbTz9Iu9g9cZhLYSIFFaXEr
Y4RpQwkWY0mg6/4MOKgoytYgx3WIGz3FMNkTVuuI7EwzRvOfgqw5klJVy6ZYLdLU9WIZHbvFFf8n
0VtHKQ8fTKEwkNLbPpvfsYMmTQhIt//qK8CxG5ZH7s5yo6mt9Pmfxpa1HCHpUb5oy6HK1umHcl5X
VFuaJzzgrO6eP7eRWyRgLICx274fmFCyQi9k2ioLN7A85+/BTx7vEEOz50yuMSMawKGuYDlawnqa
CYxh84S7/pvksBvIfaltD1IjsohukU3EAKHOHmU+NFxpmYZpOZpu2dAeIRQnrkWGTn9kryw5yfpp
qJlAbMcEC2CZYUmGtCwacdirKPWaSHUr1mSXhrPtYoAHHJDpkbMEWCy2P8QfzRckIB1J7P+L0VLu
TLBAVhdy1ePNjhI8oUu/zyyfEdewc0WwmD/DE2fgVMQtug3eellA1g9WDnZXuiXpYfk+Xw1hHapI
OPR7i6QL/6Yr8lmt73c8/sAFWJU6WsMBz+5m/CIqDfw4JJiM8Qy/wkZiTF8Rzw4Dzt4Ufo4dAl02
hPBswjBcZrZ0mQtk5s0IzgNdQ13X+v2jE2aO5FNH5iT5omc+WPr94fKFRg/7SOPBioTezCWpBQgB
yl8DJ4ub1AK4D9IGGfh0WV2bqshq96xwIkrzrckicHHXPbza/TF7zd6ZJ3aYHmEHJezUWnowKqbE
Dd2rSC8E6+1aLEgIm/BRgOYX5tdO2Z9tHe6W/lhUFAcGvt6XsAwkUkhXeDejhsHzzh77BPYaOXcK
XlxY66M1aJ/2hXx5PKP5XMBB5rbzIL+xOHlFuLsCSthjswx6dg7aseYN//vOIWoeyjY+TXUfBchF
lijJmra4ZvtQP7vygptzJGAJbm6YGaeIB0IFgTXLUxoVfw6UdzNP5rNo8rqtA4O8zDcsU1Gx0S7E
TVIPoeRGe4WdJH+aSYXwpAeCHccwROaWIw5upuKVZriSumSjxFXa2/AmsZeNL2/i5rfRDEWpT1bC
KjuWGdLXqYr2ahqFkygCcL9bXXPQUcup9AXTrI+WUMpkxEcRHTSDPlOqqz8JgkMvD4HTjOPozUYY
LIulEa0FP4EQbGQ4tWG4WWXz9RBvc8rHvcpuuOMgUlKtpXgQdrlSNqWvmiwH1WgIi+FCs2Qj8Lng
mKURILnzglvjPpfa4fhOwWPxz3rvzV8KqwfxRP4Ug3OVtR778y4odGvU3rSdLkjUDLAYUcyTokpE
YQm5Bq6ILcdCa4MsM2M2A6mDFOj2M8RYhvh1f2BuQRm/OklPJZ8TMv5lRQuh5cr0cU1i8FdFUYdH
MPhNM4kIDJr9UewqYlHRKpGty1l7GsKBLFfoUHC/StBvXaAijxpdfvznHU2B79bBofX2bxBaz0mx
2+1t30Oyz5aawNH8s5kEFa2X520RKEDN+N48fpYUTyTwlXhbKkHYVgWxUgPIVRdymzql9x3Xh8oO
O2JvNYLyKc8VybnUnYDWt9OJb8uJ/Hd5hy4hJzHyjnfMin7uwC2fky+9QBGfnZzQHrfiJt1MVPhP
V7fGvXrK637rkX0SagL/8FIejQUp2MGekh3RwnOKG9hkOGnSYuTQLhXl9NCBcWpkrXxed5fCdLWM
q5dLSxeEtxaf4rA8WFw1ytXchlWoPdJZCVQuv9ELS+0ASNmmToaHqII33layFS5h6qKVK9rCdWLQ
CMRcyxJ1c7NELs4f44E3i5XvDjrAkiCkCnB+p+Iws71aJuiY6UzeU2BGcXk0IjN/KQb45cSfpjm+
ctaNjsa7LZ7Rv4ArstLcK88iCViYRv3YpvWyBOHKgoDydZsVuHSK4f3ocTR4k9kv1TPQd1C9so32
rYxL7exWhAeikEWU57Vkf02xBfCaDzESf3Iw3OViDRa4mgxSLKUmoziIYRkHk9IJY7+RVuvdnEUV
1wK7VClXxH6s6GWw3FvR9CDx+xtnjztbJFx4gjb2HkNPZ43D+WsvwCWbhoCfZ+zjKFvW41pxHNyX
DvHAsWlJx40WzqalBTjCRp+CgrSBgaDHmaipJmd/9RmUUpSdJpkM26C7/M+9RaVl0P+mGqYcHEn8
BJrG/xHy9FlVAhdDG1+Od2Zx+pd3AeKXcgNGJQ4uAKUQG041j72kyCzWsl/d9+tCHluHkPj259Qj
xrJEHKcpqH7+sEQLNkGo12cSh0cHgl/90o56FI/BUsRYUymFfemJAhfodiAkA+4KbYUKAVlKJ9ux
eFokM9Z7foc4/F2sRuCaw/cQmkoVPZ2vRvMgpwWkCTcN80HE4Ql4xJGOqiRGuelyY0+Fr1h16MNZ
2snUFOBC+mQhqQE8ev5SWyPIHG6sfFwWz9Zhma8NiIP0mnBrG0RANVrb9COYBprggeKAGaQzWWZY
HDAtu4rVScZy9m5QKJcXMtG0EC3WEXcdzv/g0+wd6qn75lFEnW8bSKHKzJCIugXrDnHhAt1Nxm3n
bI5OzwQH78ZpQCqrK+4+SCfh1dZLlHkbaxCPBSp9+A+VD7sN8+ZUjN232K1fZt7uZAvC1sl0sXNh
OILS8HGu5uBnxs5WHyMkfB/rivL4c39JF6WYloLOXQIjZiXmFgCOlWc794IAM6vcnqE+Vr17ieUV
3Jx2qWb1rNSjlzkpkiLojlkd+ytIycjMy0ivesgpgGh8iLWwM4wXLQ+eSLZy4hKL8tvpSZZUS4QG
6Xh1fGfkYkkPurnwSxdrqnQYE0rjWm4uQJaTpUwSDMimlXBSS++HNVTT+XDuw3ESQVCs7tlRWkog
3P7gkPSbV1G/WzRdGeuAvvBa0oW/q/iotwxwYd+g0N8rkRr+ePmyM8Io7g0E5KrmxfjGTmK+NnOF
CNWa5vRNJMyxY37w5TacRVql3Xt5gWdTiX/2qVsnvBFggirTVYIZj1deffCZZDL2WQw5Smim4j4V
SxPaaLU9SjR6pZoEx/LC9Ix7PAH8r947PDdzw1yWaYMv1/x6HLzvea18c4X2Ju4BXbwPrvVpH9uM
Rn2s6Hx132Q44+pg0dqzJc9OYPBf8pNi0C2ZEImFD2zt7+6R0ycf+2nV2LR8dB0OyzrMPLbbXBtP
cGOaHSIsYjo9HibhLrfuzq4faG11VuWUyzSN8wUWTDBEjPihnjfEYNRH2U10TDlkzK4lUniDOytw
pGbcSDWxoX4QRnwcLTwoQJCTVUpEUXaQDUSj77x4ygFwdZOTcKEavwDwMhAPcTMdUemj68bmihxy
ygXPllYzyFFgOHCTW3oFmEEzC7V4CJgxHfdnIrYmSeroQLj3ASeKhItQOpGvalu8brT4QCimDbnK
AYfZ1NaO44kX9T5ShAVvOJ4gL5J+63i1eyrHm7FVKNxtLCkRR8JjnNCGDVWbRbKQa9kUUP2brpqP
+yoaQuV5N1FkgjPMPoGOC8joFBabacc66i6kF+31+D0f9Exm2pXa2Ilts3dJNwrOf8eeBVyBC+0Z
e2tG6HS6ts1uv/wApdOBc3SIYCSwkUakccqyKJY4dPLxEmIFd8tjrdjjUoPUIaJXqHX083JtBcG5
JrQw0ifeeIVniVZPDxcNB/+7AULGP0/eybsiNLDvMWlbgce0/xl/Tcp3YQFDGb+HffuVpkMcusIv
503x6/UO7mMP75DebsiXSu9B9mUx5Vs4VBvy+OHZ/MJLQihAUk/Oo6wo5Tl6/zkydxe7q5GnXe8z
PgflSejz+JjhccySlnTnr/xUz5B2ldgsghqM1eiW4miRfoG+6kaztUE36aTcZjsq/IQhR2DHukc8
Oo/48NJyZ73QZPKdH8AhYSVa98qouzmuwaeNT03QcjMw2OB/JqWpVr5v78468ifQxZzNyBarzBSx
oinfX6Gh2kvxNCN5VpL5pgj/WZv7MfrI+Opi4oQ5hTiwkDNkhvb1vtZ9gqDBCFvENdsotDvXbsCP
m/0ThShoxsAUWLmnbPUvm6gsoo05KamBFkThUBsYlAtX8W9Bl5hSrqu6IyuifvHLpm+bazr/HY9G
/SllvnRHRi7z4qA5alRw5shr3yaoJM1tJxumKQsD+stNwvxmazPOpBCGiZ76E1TjJaIFBcx84T1H
hZzSCZuhllM+1XjvHQjyqwFUdELPBhGlwKc6hOvHhh4BASXPj7tsuAMFbbouCEugF6mTOWfUPzSc
l9DiBN+RE5iUW3E6lvQYBDBz7ljlVt8F/n/3agtKR796l0Z56K8HHxj81A/URrxEinC0yZhGFbG2
Iyv1KZF3GWl1eiHjMidIUqRjQYRhOMhVZPoA+9UlJ22vnNJnRfI/AgR473+NVvwsqF6VRZC3pyfF
KhCwpsyPHNJEVLyDg5nzjLhreW4FDH0V2EHCLwQ6UcHO9p+WGzuDKp9w31SuGJv4ivZVF6rO3otS
jMtcgsNNKQhUwg6Uwl8Uu8WqjoL08oz9vImDGnFdBN06Ymel6UbrTRcnXTl/WdrTYL1bUsyBBvKk
GjfJ2ioM65IrFMqaB+vQWpmLtsbkS9l2QttR2Y/tABK/WPSN2+8HNqOWyVK1r5rw76YBSqg89LlS
I/DcSxCM0J7J1xBMtBlZ5EGZ7vrSZVeElEMMamo3YsuJ6tpEN0Dgd0+OpPwcFmy4ERVHDmSNaF8m
Bjppk9DJy7/bCAJ8bSWROsvYipnvh4xFyezi0GzTlePbuH4fiUzSwVC106VA+BmTTdZc53PRYebM
my7pV14fpGJGp29KTblnuuH0c+SfDsqgzhQ/l38okH4YZjzYTtjTFF9GhzBj2WRngwu0FCb58mC/
NhbYsvi4OM/I9HuGmj3fGJQGPvvz0iaPll3Are0qNx2zlX0Tt2DE1GXO5J4i2WOTyc4AmQLC6ma+
SAsPuHPfBn9XIBe+E8y1TQJmQIxK0eHUAlCRd6Rr8meTenwfuJPBgpd2YXMAui56tlxpI+5f96E5
W4r/u0N3oWT5C0+ciHYOpwPbNSDvUtPMyp05MBeiqnWcgf6r+YQiuhEB/friFtznFdFlxm5Tsm/O
MYqFGTAJRmmy1/YgezEsMnSw3nYxCiyi+4FLexoKaSYv51UQaV558imXWj2TaCbZ7q/Pj5yoRp+8
fiA8u/zTcHqCYJsDM8FDr2epEpxRvm17+egXeAZQ7EQOudFVFHVLPMglHqsY4dEitDMZ7Y05eKrX
YwR4hvfqbcCh7TENtqv6d2x2ZmxW+8Q3HhFPnNd5BADyT4PoNo6PFV5uZJ9HzHNCG/9+7lUFQ9eu
/auDB1BN7ygCd1wFFKiQU61wZ2QPuHJ7JSvEkILWyDHPR8QaPfZbJixFRDS0diXc0lhuz8B/2Cz8
rjzgJSvAKf/QueYJrm6E/jIogusELu7Z4SwpBvxKdpCgH8rtyNojv82G1mb3p/ACjg/xFzVyzRqC
5egiYI/CpqdvU+XbH+JSVHGhOy7T2LA2LIQ60HRq3jpuFyXiwLfC1EEnOQ3X837MBrDnlSavv1Pw
qF7+65Bco3ZCs+++AvO+IJbeQ3ViSYB7w9PCkbJdksQjzkwXk1v9fX//0bIzjZyFWTcUVPq+Fisi
2eBMLTBMCB4wKv723iWqF//IaANqwx8EHE2glAHIl4gjXL7wbkU6eU0uvzeOHhuhXpkMnW68Nb5q
BzeEumZLakESo0oYjrluf9W2yTUOsn6QpjYP51QV1CUhI70m1kD6g2QaolyelI+vfmb1OSVNRdC3
Ju3CS3rmR0zMLks6w2Zu78KRMBgt7H2Rg5/HcdSbu+G1ztJn3F9xzxZHs5TOB4/258fI6OPg+178
duY9qeunZBPrHabi8NYA9EjlnVUOv6alE/i0Prc/dY6RmAkvKj5qpRIMMSLktEie8aO3b9q8amat
PCAyyG2/p1EBdDi1FttbyIblridXlz4UYNAKBQUnp19yY9LswN3IWfG8ZLYo76zkRoSyaOvbwLqx
Fv4zBZFwtQfxvh4jnnra1nOnDS+ao2pLnp2hbd7qWzlhwk+rjMEEYxaITLVdAEFTvYfPWhie8C8/
HnFtr4x67FN3XxnyciL/CS/n7jpaJ6RwE/PAwVkgUFbMEA2FhAOasyfh2Yh0LWmHQE5hNbkrwrQz
sPIVGJfOxeJ5OTfGAKDBK9wez/tmZmFj2cMH9bwymoAKGYpJfXm7FFEoA+z/cVzDz9XRf8GqXIpg
11Dwfx1B8CbiGuzPC/9QZyswIO1UBYFSBT8SZP4cZ6+ZWF4xM3i+3+j4OPcqeBugUUl5oPFfOOO2
o/M0zFeC5iOW3EB662KCLKbYnn/VEkKCKRcqsfbiDAZr4IfYQ8jr7WfoMFX+g4kZE7gu1+TMjXPt
zaaZxaTzXe1T9ROgZbP8jimeV+QIEwnctDvC/urLxwlQ2FcA3VRvT80rP/CJ4x8PKlHsONLLeK+1
MS0nsFf+qUoCctZBbMOmHTQuGmR6nvO3POHZMAsrWQn3qPerFcnWpwNGE8uprguU9VhlBa0MCmme
sjbyO4pKPFoA7a+nqGibumRG/D46m8lwrnsW3AiOKIHXTzTDtmy44HditqPHdGzgNMYKbDzJktsk
tWOy1NYw+mWNMz11d9orPhpC4Wqluwpj3ng3xi9yuTqcQ+3CGGFQxK0bile5kg6Yo3Zgl7rGOwVx
lgmMRfVt+ktTfJeWSeetJhvodtDNO7WCCZN4Ev7mD0CVJew+R5SDEougt4noYCv853epRYXgXq0y
HLJcUVGIuk43QTWnftanToDcSzZrJlUDsetVWVYR+7RVblCULleabX6qmy0hk03lnXsQ534TURcw
MFa9ZHZ7GC1fsZnpDpspUc1hDQ4ZknouwhGj5P+brNSY5jFZDjFK20mYi/gxwqdV+iysULhgewFK
qdSkSVhKPPlsZtLuMar3APeTcPznxtn2uc2ef6LSGWYfw2ErguSJ/9Ibs+cI3d5BG9pKdR+5M4hu
19rzXgD2huyBwfiF9/qD8JM26F/IFPCrQccEGloFKR/lFFTAWxh9+91OqT4MthoOazIUSDw6Txwu
U9FYwss6jvqDzyOTmKTGWsD2lgd6JFhEfCtWKDLlW23Wjb3eakJhQwf1bFvPbLLySnKa9bnu2Kv3
0VytxNUZf+L2k6q5OxCfaeQeR5+mS6mTkqOBxbr0x0y5EMcQA3MtyuqS86LHHqKtp+V7xfoc3rEP
/VKaCEwdmjjGcZf4Aw92NgxyeOkSXX3wjlp9iuu9pXRBKs1mnIogyCW7uTrw5Od6jbXSyfBVYsZN
ejPe2Dt31ylLpkLb75yL2xojhinFkvVBZ/jbXgGoDo14eStXARhvCi5/dZk9ujTi3U4mWEJjfIdI
aNRVswzwrGLaTM9dt+edj5/oiBcQpfZTDvRwfpQfsHXIfRrV80bBcB5eZ19hk7KerGCuIE9fWvtS
ralsPiqaApsWXuIHgy+ziyCa5ahyfhCbFcB8EdEpilvMBj7gYwozY4hjvnBazMYUAkcNmhNOewRG
4pLlDpYn7wQzMnD/DLAHCxYnRYvYzzQGmR3Q69/8ACZgQq0Nuy2VVXVxPE2RxBheQWbdswOtRTlT
MLA2RjjPpSCGnXHNoZQvBfv96Yvt1n/+4hnrxQxs7LA8nKBT2ZvSCSaEGjuTWmyS36gdrTSf1nao
5cXtcOX0y73UCZkzjImwIOFg20FiMA8vxnXieppkB0Yq5vamBftkJ12RKG5QCVbCgzkhoEuDB7dd
N+TvtQzPDYCOTDeJctkQ2sMgxwxzl0V63fudQTK8md734rW81VF6Fh3CHmyNUiimLHGK0CtI0IoG
4nKl68BG1e6S2r47CWXg7tN2nPPLvhHiz9nK8fNLAQtKAJd/7RBfauqtMmv28a6+dYy/PKKse6+w
Javb83dtzsYvEoLb/+0I3S79cvgzUcWJj5TRm+4ipkTIOSPI9a+okWieynVsd5ZgKjCUk6iRo5zQ
CjvDMFZATvYirkmgHn+nUb1MfspF66GPos2lZFHHSq6cLOGDd+kC7FYtAMApYBfwMlbVvBomNrXI
C0fmump+HAz4iSjA5vYI03m7vEmujRYVdg6b1CanWzWNCEkEZlikqK+aQYjkcUYJMdFGdQse+C93
MhLG27sCUvOpD8u1LTPCAV1XMIYTyL9TCCrYuPdYyO8ckdfeW+LTwGm3jDnLeJxesndy2ZEyJP6B
Ufm8QsUMLcDyFhWtjiWkThY3FOXlXIwT5Ti9fyLH3T6y22pDnL+kX7pTE82QmSE1anE60+ud2kXp
XD2dSE4TCjl9+W9qUGh88bkm9SghgxqKzpsZ1qWEkXK9mPvgi7fkp2KKJWbT+raNeod+9mm4rsEG
VltYsbFisz2NjY7CQB9TzNseqzwVSykmZFB13HJ19UbBsBnp5mbXgbKKCOW3dacekOzIegaEFaR6
ZVNr9VAero0zF2cWk4XrJorvYCH/35L0NvB/IvWhMjltGpKuj7jLxubWfEkBeBchddFkNXiJa9Kj
bfYgbD0oWTi5nxpF3bbmExtkGBQZuXHi7qd6xEk0BK8Ak2C/dfnis1kRWnMPFHUhrKuTXUTWj7GS
o9WMlLJ7In2EeBNFQQ29pVLUGAoVFlyKjGd64UOjQjJ/ZIrvRaLmB7YlxgpJzrsLnUphRyYokYYD
5aH1XBm/DcDKn+a6gT5aF5Y9HYfEMfW7rAbxx8+hL4mJIeCQJIUUp5A31Q7FHaSI76y3DOmjQ8mR
Q83t2S48zc1nNO1UQapSvkYjR3w+JhZiexkC268ts2iK2yeM0inSEIVJ4iTF+8tywa7WmVFgwkaT
sHIqC3udlksI2e5n8wwdrfTKs2V/Q/dbZNVDM+oKTYBFkvS+g8Ce9Gem4KhP6KxFJ978PrL8irTi
SFHd07s2gZYZnUHlOONo2EGHySnWIgVkSmLx9FpkuAPSKfo8dA5Ucpc9+0NYpwXXHM1zTHy9KZz/
ZTnAiZp7UYcEmb3O30FRvXnAh7lTKIm9vevzD43NRDIvA4ihEIqfQmVCtLDhgoG3ZUkBVTEJHE/b
U1o6KM2OXU+x9rwJmyDO24ysCTrDkszPRnidoBj0MpWCcEkTUQTHJxjaHzImpz4ljGQw6mKTO+B+
Q5H4vDdcFOVKcUx23iDPMGuf0imoxHsnC91qTlYf7tfrKQXRzOrC/6iBCyw+8PkuVBBAKL+J3vai
Xtf/UXsg0r8v3mcwPrMTY9Cu1p6rqRkOlu6aNI3eq35hVBvt18jBr8cT5J6FZk5Axo/r0xqHh2vH
mx8bmbeOrKjYPijl9SwAYAjiehwpmBLh8dLwWsH4KqxTY2aLbA5GFwmRxKnBSY/kLUr+lk6ViRTc
tECQrrQN4ncKKDlQ3CrNA0OwH0FyVqNhFEIX2VWtHXw22l7kDXsDZP43VfJPojylsEuvf+XHhzNb
wVbGg46pXlpTCSQpPcTXQlY/IZ66wtBdD8VQgZYOF3vbmdqlx8/GLmsIFjDGi4Mj+wwb2vmONxUj
+MfIKEVbn4zj+2x1jUSMMdrDMrU+x7PoZGCZgi/Pa6pOafygKSpehFdFwux1FB4XTWmfCyyvjzba
Gmg+krKD+MdmGzbVzpZg0FNg1rzPnNhLrBxW420lxuZyfOEWNDarM29yuyxxDDpIn7pV0gV+3i5j
elVSVGKC3oK73sS/nkyIK4p3t3LQmqiFjxlPEbhE7PzSjs6bsJYAx607soNUGSpyPsFtebB3hos/
g/oeLupJMSoQLOFgkpSZvXvz7LOJHjE51us6PCPYEtEIk0GnYE7cW1TQW+m+tOGMp0VOUDpMwgGF
VuTxVB3Wl0d1h/yZrs96jg9DvEKLIDQG7MsbEcP4TXzgLB2WnF46InkN46l3H+9xOjnW2j2DC194
DutCawXvuhWqCDwd7Md+GD7PPfonwOGeU77mY8no23YxDa0CsxLVPMITBgB+gw1muljoG1SfWU6a
lwx/plCMbCHHi2coeFAaDmgM+Ka2munInD8vx27ZNJ4jOMLINRoExuqCoJfKv4zvSyvVt2DxGiF4
FcAG5TOa8MD4oyzZ0b4NqWmzVMI53Sl9l11S1DYuOFjYLFdJfDoBrI3/tu44X84zC24Ms6olEhR/
qoAdv+gXsD7mc6WUEtEenhvlb7/t5njtTNPJSUAPAePaYYBKcv3pfpaHXqXusUklJHRfObgHxp9y
Uv+xgmEE1zYKwsx7kjQcvpVpxrmLUZQoxV3t36oP2wDEXkVJ/TX0LyfkdyRt224PB8m6EtBjFwsq
NETj6KVBoLS+CO3+bWttYrkBWIOSzy/nAfzk4gbyv71LhRo5GP+TY/OmAZkWR7dTp7Avnm+ExkHl
uxmchMCO8ecyuu8i0+ScT/M8aNjrO9SeGhFz2ipVs0KQvhX7B8JGST62sgYrJVEGa+B7/XSH5xKN
JrtpLU3bkLK1bvtv8QtWby79B4ZdAwdORtz3zMhwUQlusbGaA9odEqmHPQWkfMOUpUdCw2nHSAJU
Zq6X9/7nGg/aiFBuBJLKZmL3FIITcSpftereqVNOjYkEjHB3WIPMJAbLoWDR9xFyeOAdj2sHAK6t
rTzAwe0LhauM4CvxscLdJX98J0bSKRGTC44tqrwraViPJu2wg7oekNgOcmV0dZXNhhvLNrLLNNue
seNuPfI33KIQ/HfzoSQbNm3qJsYqMJzZc5S4qYvikgMvhVttGiDrJIoJaA6MPq+PctvcPrMquXI8
aX914/zuRj9hjwNFDJMcBdkNBLWx+4HztsOLLg8M61O0t5M+fZifQ0kQO5516mNgl8UMql+EKTQT
dsd+1sGpBMEChshJedQ5/KFjm9srWfMCX/MSO1xD6UdIRsykq9HmIV9Nb6EPbeGm8aqgmgyL7a9/
2NIhtbrwrICWNvDJzyjcLhcS3TMNjpnIjfJQXI/T+0nvxAYdwbQl5Y/qYSaisIN/fPPLF2/QzdIf
KbbnWMjPi+HONBcN6EkWBoQKNF3OnbMfOVTUDEKD3CrLiKOqeMzMOFQ5b1jtscOmrT0XaDWlDpuf
05A7SL2W3Vo/x0kGWVIoB6d/X8DkndANdl2fNHvEI6FQGNWEzyQm+JlhTPxSyHaber1eF5FpeF+H
rrscBBegFB1QsH0RUFUOj2YB6ZYsMAXznIse4wVYYrjXxrsj1gg4c7FuR10zRIkBjxhm/tebRA7b
i1pK2vsehaUnXvLCiK159lSuj0e7leOzjhR9ojKoXsAPWBFPzAkxw0dPmZ4+kDW1OcA46sVoc8+V
7d/dV9I6RQrj7GqWVqiH4T4N41lZN6/mijDSnnvWN5xTjLX/gOx0UhNbpLWkHPyQj8OJZOUwEq0v
I36NrQsMFXEWYER9CFtUvBQzx/6QoY37QttlryUsjobd6f2OX1cCe6F+Fvcv9FtGZZ+AHtxmoDbf
g2eva3Pp2ZZAEaMEour5TvqmUzzaz3m8O+xkMJt8kDowMqvK+5bwm13cmDsUg3upp1O73WXLcFG/
6gbyNvHNtiFNgaYWAMQR68UBnuKw9oCSUQ7CKO4UPUGm/Rj9sQgPCp1NtPgSeJTlWzXsxDTtEpCu
gy70/TRYz+hEXtcM1kcoAooksqhHQ5q+EpS+HlLbS5WfzTVWInJlSd2oIek3wezI9E0cKMpDIDff
TgFcHdqkSjo18pmr/vSY0qXH+bESHcml9NlxUhtDelY0FSKfDAZh32EbzHUiiKD9Dg6jr+z54sya
1mA2lpTe1uwpEvf2cniNbEpSjs6cCoCTNt5pZbfW0l5LgDmBOSmD3HnybPUTPLVfNuXAvq3erQ9W
gSPYBTBHyjraTi8vz0Sg8OTX6SbVrkjCP3jry0G0thkIQVaRd+7MzsYBTx8M6E/87rvmURGLuKCm
4aUdDKEGFQ/LCd6MUZsx1cRWNXZhSCXAtjuwm2h7l0nTVWQQolGAwzNYj2WeK2ERCwR9UvfzOR1O
zd2qv7fAkMmMqMor1sIH26/fxyaU9k2gpC+TTTuyOs0Q3WriQS2cdzuCKz/I9EIkB3neLMVMDQd8
GCYmnquaohnWMXiSrm5djnK3qT+P39RzI2wDeBZhHLONWFIUG9mT2xjTcO21iaus3DBIBtgdxfkC
7n361GTpv3nHar/dLACu/QIVIDDJ9v35FRHpEiQhcc1agvPaf1LqE0kkf92j+VBTb4jplpO9kVqm
FzP7ihp3Zv5jomq6HiQSadH7mitvRJNAHJAgyGSyrt9SqfTnd8QFEEnhX5Ixk0QLuGhLFMl0zPv8
eYN0pH1fuqjwfzAlimafakY7bbxoMy3p3NrnDX1bRvKlKKH8/lyAtsTSM5/5gx9g/Q5vxJiijjSd
bbJD5J02PxIu+gFLkodl68aSgiJWSBKwWdjnKZNmCJ9m5g8/rpf2Vb0eKRQ2mPRt0QFgPT0pv9h5
7o1vFZLoHFizYWlD/Ib6NsYyncbVCff+PxXICnIuIsjWJym+/bD5c5vdn02sLhdebXpDqaQdC67U
zc+Bx/dBE0wPc4+jjOjxqzIa3CbmYE8FyqcW39fqighzCqS8ucNj2ViZMhNIaDEVd0RNKWPlRTeX
ZpGeaUby2KiPHZcaAVjIGgSjKHEII+U6zYAX8FRspePpGHCrUK1KQo0BbsrrH3YrDpmEHzAIPr7M
ouSef/0oZF0eg1rD2dT0tGWLJSm6ozyaOG1OtYmxeQxxqChBKkHBIZF62X2jp32l9oPUGnx21AiE
4K0D91mCcJvo4JlxYjBcgeURSPBhS9CEPgQNKB0s/LKwWIjQEol0jSbg2VrDr3qGlD3Uq9JeGjC1
1B+aoXBRQKM6C63YSS+2NYDGANnxGZZjFWeDvJQ3uZMYrYne2Tm4I7l0474UnaUUV0BRshGRQjRi
Tm6la85YRGHZRXD3Y1FmUhvMgGPS+tsWWl091i4VXTLHsoTl9Exl/O7eNGhj22OE9ytp7E/ohz+E
f+Zq8I+950UTmRJkpwHNU9Tzed7B3ZlUrZ1uYT2X6sodtQvu5A51q7dlJvNeHUjuAhpfF/90E9UJ
oKd6ZIbOWsKspItW7l9fl+F4+3/njte91mad9MT62ogTV/X8+KmHEu5rcxp/f4zbJRU0KdacjKke
jwAjEgTNhcTz4/r7VyYOZgsGWantVbTIpwkf2AE2LDh/Rc35vXarTrapc4uwJG4i+AupabYPsvZc
ZqJfIFkoqwu7SZzfbrlC9iZyPLvZj04AfQFYdaUZkhBoZte7Xp/isfyZeZzUvwLhgzR8A3loWfB8
YY00irqXUHyEOBWNMHWlvVsui5H+gdfso5B0pPwqjtdSTAnZ4Ll8w3Nqvk4Magv/IxrqLQsJjyvu
XZBx5J1s4PmeBDGZ5P3DRER6UP15RJIcSqFAKKCPmeFbUukfutdIs0vKUlvHMIav8UTBhFPMZ/N1
La4hCzBENMN8Js0zmwkACNKDGSQ6e+lYFPM3FTf1IJjYtEgKqLm4mFtONvPL4TF3ESSmEOmiA2zi
5JJcxx6lHF378aZPxTwpLr3aqDsW6x6VXiB1n58evuxzrOAQXFgvfcr+Y3IQuRjXIk6YLsZbrIEY
bHUHRhIOTvl55oavw6is1bz7Z9nYTWeTw6O4Juc70I4B6TC7nDmQVo1Wvftghz4FGPbls12Lk+ej
QjYIZwNi6wzOBqbsoWpvF1XdreIC0XL6lJxQd8sybf121Nt0cjA28Vfe+d2MZgTzOAFGOkOQxzs1
C3+T7wFBgZnx9aLMoM1J1XgF7ocRmOpnq6DA9s9ycsbI7wjnTGp1aLCeOePT4/kohqj5NHR7gL5H
OO8nltyynOHMJiEFwmxgTY5G7fgTMQtbZwxvRQ8uGljVcy8VaD4AqHQ+YWYl+9t49jK9si/MGV7K
N+4TZQ1ZFvb04LWjwx3W6UgLOihMUiNFSgauEK5wxqIhvIVSGLL0LlUN8koDFz/5CQXGWsOFkd0P
PHoGxFuz3u7aGQEC24+lvPObBKLdlm8k1TpCARFEkZBdDQ/wDosw9iAPuKP8dLl1ejHKXgnqKyzz
v9gjJ8zu4QyPfIH4lFQ1tUfpHBc0Rfq+m2O0f/s+cBi7aRHaHQ/6USsTLH/4xTBj9PnENUvsIhoZ
6uQkUZxrK709Rwh8LLnWJcYhW0A+dd3nlmCFXyxaYngEFHbii41J6lJNDKawBoHeiPuwus1VtfUv
5p9X8BM91LaTdav8NhSyZ6gvHR2cLq1PzPPjzddrN4ELYQ760+6MRAJdyWOHo7rXjVO8DfDiILNg
xPE7jlxP3+hzGpGzAI3gKvYfpa3LJJMHR4vpHH6IpYENKGPepU3fdTzs9BIOpyTlTYZUpPlG2fjo
GS39pZ3QuOtyt8S0FmjOorh6eDkV32LyuFGwLwqm3+PwihxpGLa1YM9yXMhwxc/04seiUGzVvsgM
NYUwSQtERqX0lvUOoUIAzEwaH23RljKp2sC3Bie83liAxwSDfoOaXZbhETgTwUaAnke8v0w7Lh2B
a+dKK3uygR29800HE+GjuCb9z3zotBU/pT089wOmCPnliS+SpgLHqxQHI9HGkEVEW7F5j2tZ6dQx
/GWNLxEOop34EMQ8BkFAuOqwgTQwyVRRiUwOw9XCYIzo8lVq6lMA/tRcJvzcqEyZ4rA20sa3pspZ
a2Gn4g0mtYi6oVynA/jeap2z91DDdb7zlVR3rdw60fRnKcY5XOKt7zMbVCtlkFXWG/tOuSCnLbWu
wTSHYQQqxuhVFz4krvsjTqwbdJ7EmY9qJ/sIRz2HoKDLsItmZ1wK9asGhdjleqoGsWAM29q+218d
aR73feSzGvh6gI3y9YCqEnt2BmQyktcrj3mzY2rD4QUh9f/OQmmvNwrQRZha6x6cbU0TYjNzB4Ob
YiuGK7J7SBr4tioIIBP07XSF5SouGPosZ63Z2y1xT9BC0XqYyAvOaVH0YaDV+e8l5T9qYcLLZUx2
VEUdkWCnyVYRjONQYM+HyG8ducaju9kSJD3WsfYYfA8FLSMXpYij6AdGiu5j9/rRwv6E8BMyteUR
OGLsyODkz626Nozr9oud8hgE3PESTAm9a0cSEXc31SvxmrDNo0YaPnXABrXNSnuBM4WUBT9rGN6Q
rU9rhf1ncdPxGNRr19JUyZO9fVXLD1FLCZS7R6FjUmO2UynFNiDrFGdnP0iwR+bNnbFBmcqlDcDa
oD/5JPUGgASq6ZZQbTzfWzHl2M7YtnlNhJhvWKTPw2DKKxVmVcewUoaaFGxzfTJuPaMn6FRAeKCN
rd08fTtM81PGzRL0dpLRzybh4qb8LAtNk4UregScFRUWKsAr75g9u+UBPYKL88Sk7y4cyjwdAw+5
t+fAqfdk53fWT2BtD7/yiiD6y+tGd6moauWDevrI72zM/Sa99hD4fN9YMa8uhT/DKH/eJrb66rXv
2i1VaHZhiuleskHzt90YbDBwomKUErVfEQ3mRBQUOFpf6TsR+RwQC1+0q8IfSQPbteR8fN6ZnYVI
6yw8GDKvmLM0UgSD2sTv/r0Kbf+ZDeAQn4J7/I9ruG309WYhvrMXwwzewn8xAHJpitE6czL12twf
7lZ1Fcm3ImnNRxY97cfKXIh0YUEaKu9vUCNynPRdDSAMjSBPCs1w+2zVAEIXQd2Qe0xWMuqtka7n
tzY0eiKhNLHGHRMTWQqwYWW1DnM60MKoV2k3L5hRHth9IJd1OSLIy6/pNQFhBqipe/UqG50Si0vB
ejjUaKLYVuclfPxKkmN13lEgEBxRUpXFtV1eGo/T08zWtOgx6TvLvgQfheYbrl96FmTeo6OLe3aC
CbGHKpXtj77Wnq4HmZOcGakk3QBe/TR/hEYFkJun8l/W5EMaMc4XWL1JVWiVPYmPviYAV9NOrAU7
sEKCHN4q748ZM7QWrVW1SBhwrYY4d20y6qEwz/3iB0Z3dK56qyuqIb/3ZGJukd/+pp0r4TVjYTH1
lsgfmgirj908fympsGcwM8MdiN5RLMOxjG3g0lWD2/SmUCwJzByeQ7ZmGxRNUSFx4f6mz7vmHuH/
Rx2sH2cX2FJ9HZTVMOFUIdSF0rU1vg3HmAkpR4hXCELBwGkA/EmzufgV22knUwDOXY3+albmd4H7
/NEkGNGUCTMVZtkczv8D9jsO2lFB8PUMnYiuE7erygrHFNMod79fLMAgLjiEsb02elA/RZZjqXGs
EiJsvQZXerAQ7z5WV+08+cVnz5rqDyk73PFDl96d9hLJ4qovhhbcM0Ni1jTDShQGg5NjyvXdi3RQ
CnvoW5bdQ2HMRp/y8u7u1ajCqGNHH9BkLHH8Dn2gVuhl/sgME2VZDk8I/6Km3dsvaZqoyuRk9j6+
ooNEIM+wgGtdIfv/RwrszXUEr+fAng2F2tzfo/TkKoEo3TWoifJOheNMwMgCGlHF0JUBAS8LH8hz
rZARKfmrUk++Ynnqa9XnwVoiDmz7IDpKphVoe5RwgV3Wx/mqE/6p3tR7kldcqWw2hgn5dA7a0AGY
QofmorZPmVsXNsrGG8y26Dj/JUmmZJcxgHWjI9irbpKbSDMLgY+cMKeVRxx996qEzcMHzEPzfTnc
SkGQOP0WprMFprn8NeQtpCrH2OeYOhAcnkEIZkM0L9qfDJ1riOVV/PiQHZQLtvJZVfgyo33acHZk
QVTzvr9pVJHOFW6e0RrarlUjSeST/7z2bACNrCGcHn0tNld6zoxFPm9NoD8S5G9TC32Hxqv4XBai
Ue+rrF4n9SR604MMx82QC07tL+J8A+P6mm5j/ZgYWo4tw2Bw4keI1AW7Zu29exWaioHSgUeTpOrK
+LydRatgVCAkStMR/OF7avCDYF6hE/DLV+AeeJ8m4tduQMmKV1sz++dt/xeG7gQFVuN/F9mex4Y2
Sh9jWu0trCzrYlJqcedW/RiAaxJ8axva9uAXPUn0Nlpm4gr+Q3qRt3pwZXD+6SD0daOnGdYAHZba
06vhtF1ZytrDhmO4Fkp/kcqnDQSocH3oR7UyuUc2YvTWB3GLQmT+7AOw2ERd7fdSw9KysvNdgoJN
Epfth9d+VYTsuwwASWH8b4yR6F7cbLG46+AJ6BZEyXxuOSciCouH2Bzlba3ATCRj/LZ9E4zA9Ir6
DvDTTJmLxJBakZLKvFHMv6csfztlkt5k60xDA5dHdmgsQLwnzwdkmwmlbw+MJ0KqfH4tENoTo5ev
Ast5hx2gLBQxuxqimKFcgpurnEcdo+sSTNWZrEqaVwI38jziPhwOQQjrqwhM/zy1IGahYxc9hhyf
Bfqj2MwrvwyCF7zNCzsvEmtJV7kMvHJFxK9bdNex4YS6Z8IAuNyRPPx/la6GDCuZuCwM6V8oUdLa
3jDaLt82JEF+WdGHbu3lbfoIsxQK258D6jKplABeSRb0eLE4pShIYuDWOYved197/oAN61659WaI
LVW3hkkc1jS4BRmmEJjQt2KDSUfxx3wnjt6EQKpXpZuSGmarSbAC2e0IvVYGzwfV/7pnxFMnsdiA
7sJBb5C7HyvES6Ebupt5O7WHnto7obT9aNEP9FDG1zexxua6XZ/6OTa0xpL4QFPB1YWqwwgY9e7D
e56cRy1vaJqb3oaWtWxedMtH5o78NIKmrW7nZRZmM3oxzZVwH0w+d22V1+TLsgxdPSSk61jl3Pnq
mHSJYPIqo6Yxsib53YYd+MrItGmPjnjoDN+KYY4KgVMjrCR5nyHhbtTlCOXLwtYuxP7ok/LmRNTl
FLLC2Fdq8DN3V69JnL+/orj9e15ydTOW3dIS/l2VCszbHKiSuAMo+TP3b+rWJre6hBSeqBRCOkNj
k/GyZx7X/Dy2FJUjHVKzfFKLChs42Pxrvg71zOJKpeOTc43G6bg226X1l4jqCoPkqTp0J7QkCdnZ
CM83uH5YWrOTqZRY/UvZqFTbvOTc8uRjHWujxiLI5rUVgn7iCIo+WMV7EoMTQCORxpUYHkVxSUl+
EUWL++ocvUdGgMOcVadIbR+pcByntJq7RcezJclxbtzDQk7BoImoBgjKac3xqgfc9PgSdU+cgYKS
Sm4RIHyLA/o33Ob5+gdAYEeOJqJmyfdKcH8Q0vmdTzgSpk2Qa6qhcfJOSM8s9HcjdxpgV6qyk4J4
bgjxqfKI3IXAOR+oSlL6pvUbKN4v5Rzoo390bfZTfspEiDKbQJAMjNUzY1lqCr5FN+0I6AgmTXNk
XbLKZrOPZ1cV6zjphIQXE+ccb4tVWdZPG30XNSgcL4LrGHKhe1TjyMaVqNI+bPAF/fVBZgg9F0Hp
yDzASs47q/P/B+TsEZXS8sR4IRVzzZ9/5P63wgZb0fv+uZMlMOE1lfqiDD92qzumxwCs+RhEVnGN
x0WICCgm6uY6FkUmbiSwJ3OAqe7DDt2VzcSasDVmjMcfjy6Jo1Fy9CRjKWneG2fWnwgTjNKX89Z5
Dg1BIJB7GDwPdlfBbinGN4V0sVkWzkPhISeyrtJ5/jaIPLTk8g3aeN2pvEyI2sFkAUYeeLb25Pez
4aWHsEwmUvRgodIXtHJhF8GtSS33ytABfGUpU7mtBiPbRXamt3XT0IPDM/tYc6xGa9cVH7U/0I44
5HCAKVVCsvcal9IJvzBsCzMHEd8lqHjOChnStwU9/a0/+7zeG5TwGi2pPfMlZ7bi4q3gcAs+Bf3c
ocRmzitbLo5/dj7RgwBXdHlwb5hb66dH7ZTluyjoYlMGmlAWyy3f4bs9qUwNWxwf5+b9Uar4c5yn
1GPZS3MDf7pjiuFc3gqtOuRYjTIi8B+tfYG9CvaCiMdSxNUAUm+CGjhn671+VvwnU6qJ1hS5G81n
eu0BJJFa+JVw2kBDA4Rhc06Pmg03jpxINdqqDmWHFwi0/7pvNq8xbjgTG/wUvnScGUFgGr5OTBDS
QWQHZ3jIAS3CEMW/mCyUXXVJncjWoumHw9IloZn+S5h9Eonel15aF13j4ic2kqSwLgsItBa7JTcP
1nx3NtFdPdyrIGvyvGztUxTYvxCpKNOG3lFo5ufz2Z6BHKshazscN2ZS/N8LKbRk5LQRQhZqN+dl
bfUy50OUntKc3Rg+IM0nGeAX0kSA+6HMz+mt+s6dKWJUaFLZh3UzgebGuqGyIYjfsIkTptCPn2yW
q64Ys4jSyY94sWeY8dQhLGjkeFEDemvFxRDoCTGOm03F86VkNtmhss3Aask8lI08Uf7B5u2+xKxt
Znx+z9e42yA7RhfSsKHgdntDTmG+xZhtB/SRLd4HD4J1/WMty+qsN3iJDAkXQZLFOgbIQxWAKMK3
XRqTLOPANWmUZGzD8VDM5TxMlGZBkcZfnVxQfipeVXLQqszr+CQ1X8kY3EuYF9OL/lcEPVExffnr
Kg/lgCZv11I+rllqgZbEwj3+gYCNqv+mWTnded+3K0cO96CGADLMSr7U3LSLugf7UzVvFk6jGe/N
C0XaX5zaNkn9TRL88PR/vjz8ieF2MHtZJueik4oy+KL5L4mlcJnCLHSvXE7XTj87NbpnhUoBrNqh
U+BkcIZkyLupYO91sh85MGJusH+t1SXI6602T/Bw1SU7VSTvl+YQSVsZws4sMUayRO5skm9on/pn
5jgQhmT/UpApanbc3K/Fej+FiIpxyytYeXqAFuf76DKOg5m+kLcGybLFMt7rZNtmDuAUqzBJvxCm
aidyYJsDB+qs8aht7giQ4wkXGUlvtLt42ass7ZhrPiWD+15JpAAN3g3GO254RM+hj59jesbYFdhP
bFlovdhMPwLuAwY2na7qANbMT48fZpMC6GxfbzKFV6/LjZhUIqCWMqJT5dvXq2oiE/tJQbWdMWbx
ktM1Uzs/w0ZZqPsP6zQ8tHFsefQjeUzsaIL0yWE0q4KFKKW/bVz4O47Qv8d26ugjOd9j7wZBcDlz
2/X6/Plw6jwDHHwTLbTauChJJyL6X2NfCaj1ut4Qi5D8IcTL7lLYdYHpJ8cT/DlxcOFQ4bmAJvc0
NUtzRzwY2R7y4vMNl0jx6g+W88s9Le9b5/RIeWOb9nSpO6RZSKzN2k5XE0h5zDTgqWhQq7wigzzU
oQ9TVjuUSqSgCynutnOIzWrRuhy8RIOxb+AXHTifn6OrvwG3BPD4bwoTMnxBCFidEF7i8BzFJfyj
PmXb8FM3BbqhvuPypYMyV5QDeUDaHv4e9ZxTdo52GF76TNanonQx4wWyVFFKLzkNXceutT659r2p
WvUEHcKb4CVKmQKmdyuXy6270Yc8x9IehrLBI+TGgKMYbxj6L1cknEpA56UUGYz7Yhyo/mDlLDo4
XW0pmG+BxCI6dj/kQc63bSIJcFPD1WgDbqEfaOGMCh1iliK/3bajOW9Aboq2FlhEyyShLcdxRIr9
JYaA3etKJ5rL9Ku7gD38ihildTbJyfgJsT173Mk4qf27iazWPc19vvtSA4qQ62kywYfAF02RDeKE
S4hFmM56w3AEN1N1HuqUv/ABc/w90GotacThMDttltwNCszZj7c/Ctm4fDrtv2CTTQpzVcvBO1CB
VO1EVOlTKVDbc5AHIzPb12/Tka5GvufBuk6YR+WQMttIH1eTyYmaNK/4Tm1MWHKOhp7Hg1Bj/owE
SkoQLIreQ6O14/Ya/rp0Yx9gnR+SAs8MM5xKiIZ1Fx4seQyjqWYbUNblMNj865YkC4bjoO8yFshP
vfetN5t1UTJweiEuHk0aO04ZtuWwLmk4ugNgxd2Dl9mcMFDq5Fulv3s2TW+cI3DXGtlvBzm6FtF5
XckneVBevf/5bBKJ0u+Nyd4aq3PyShB08eaRTBa+lOWp0gQk0p8SJR6uBegKLSPOh1AInIpvoEtH
BdHNBWN+OfVNnMw6J9aushVOR6aqdDhPwrizCQLW+5g2N4wOMk8VDAry+9XB7NafGoxG1pmYUNCB
8919eIQmqyf3dW67xq66uiGQWZ2opQHE6LJtmwGNEJWrnmqaO5dwoGmFGlTwWDeVxonSHoPmvTag
3ssLDj2/Jn3JiSYQAK5RYYg1MWw/PQrGAc8GwG0jvhL4/lZrKbojAGFtC9FxpWveWo4gb9T5GfGY
BIdbZYUqu+88llBDej6hO8ffeIWKKEH9/5O9zidD7ZMxapM36uetoGXVhff1yenjzRNw4Z/10bG5
PZIJO2dwHlg50cGlhxNHwXHdK8M3rNDw46RtS2lqCW0I2PpQEf2eiFqU+FmFpJnrPgAAuwTcLzYI
pW/BSsldjLs6Kh94ZCm1gWpa8fTzjPtRG6PqcFlrssU6qOfa1BXS7MgjWV+ScXdE7Ad7Es4WfskG
1ubFUgplnJmRhZOsYI+E72qO/X7hgGBKXf8lxWaZbNYiYiioIunx/ErE0baiq2WGqUmRZIhOw8TA
rXd2xsJ73fTWZJGj/26NLmdvCX6UIPqQ5vqyrkFCrmJMJq7ybde38FHBOcw3Mtw0+bdr7xYWyK2l
/A1PbJxmg1C02wvQa0TB7YyU+Gb8WKdXGF2ubv1Sorie9HJot6US5ddWghrQqweixBtsequ5Cx24
xvdX7aHGAze/NceeG+5nU3a6jbeE2xvShPecY6wWk9tOUyKV8z79iHP9Y+lsDItKO5CAzjor2Sy6
mT8orqWca98hvB51iXdlrv+jvizb0bY2MZqEQ+Ygg8hSHBIrmfFv89xxeVkdubIYkUZqWHW4cjaq
ZNCuP3EsVYJXyrFSSsB3fIG2mRIbLiyF39pbpweZZXYgbXI/Bfj/Et+IcA9IlwLZ7eaO5GVhXPB/
GcFtbo5RmGty0GEQ5fcLOshZOJRRzYxAVtzkq3xaKykcpTWUXY+EX6KfPfdCvAY6RwP+TKELWpu+
Hed1ZTDDHk8suLkJ2VvWl1tMe/xLo9wQ5n14aUDVepx4PUrT/C5+5hJSVhClHQitUIPL3tLVoGMM
a1H5p0O+nEYyrifnNxq57ErbhFjTxW1BMtgOE8dRFqclw+G9AqB1fL/5s3bdFqhIILwlFywpDRcC
xUwPrsNDgw0MQmRNV8P3hINJofJ7woUsXWaBTlqJGZ5buRhwZrmw3N5mtWiNWVxflLiL2zirSGAW
Iw+SewPgfFtnWyh/N3tkEykGw1up1DnjmcHUk520NAr5CcJn1Ps2m6VLwuvOV+Y7UdPFSe8vOPJ9
EVL6Gy1bnYqjIorYL67JlWjsHnS3D/0f3b2bxX986AyjtbyKL0xPLvkh9Zx3ONakQeI7MQlBBgCM
fAsSLf3VEU+Pr2mJB+NOySh41UaCvvzjucjYUTktxJCfhLfU/arLR/F2vu+RlqdRfstwTymhNEuz
16siW5eFymsrr0ZVK3uTAgug9Needo74M0H0We4sW9A86wi0NflCilt/jkmve0oyymzRkC0FPtI2
X2SUZv9r2bYTXGnxs4VfZ7hCnT44DAsV0OU6lfqMAIKuAACCscQTUzJOzVyYAyWkGwupXckuJhY6
6FOFqIN1iDjjVXrWI+okZtH3042u5UaIVwQqYBvhgCNSLEHF1ZbgAhHjaThIZxbe5mstb8PTQa9u
ntkTuh8US5yI+K6824zgPagJfR+JGsQRgSISytuTePklUv8YkCLiUjK7XL59X7d23+jZ6cdSHY45
jcofYYa1HXp3Cw+VVuITC/0QUtLNfKRX7XZrmc8NqkEeyauMkag+1ScOnM29Dvnp/mHvH6cWpYQd
OI4/29uNmsDVAxucksCjZ8q6y2I+Z/6KVLDw5JLbVETR7BqnCz0iLcz1Z+DK5m8QXHN/MEAMDZKl
S1Kg25ZJ66NffMTN+5j1J6BVOS+pSMUVWsC9oLuUDi2r8iW+MacogB+X1wb3Dwl5IHNQ0fHdvtUt
ZSdS/WefVi5kDrFlb5jx1WhpoLlTkmBnMU/NHBG04hu2O5CUMgsPkc2YFN5+x6m/sJuagiOuovew
7DuyEkP+fcKXrEjanyN83V0Va5gLHtvG2l275P1VLl7c+NCzKdC1W1UhPhxJ3WW01ChQH/uTmjbi
yrZaO6bo5iqFxpCjlyOh1CvrLK4ExZRIh1uC4T6ZUMojhFNKAXUvKi3vlj4VXiZk2OX9A2If+QDc
klvUdY8QA154fxo6ju3loJLhs2MAC3ZzMX5p3H8xEsCmk7M5Hr6PQjJpxvr1ZrmZz9STlDy2mn5R
bzI9VhqZ3V5E/UonSu/f5SsbGDqx7ZWa2T8HYd40SpJ2zxG/A31NmPigxrGexYipkSsJAO2Kvo/v
a3RsUtqS0JPFK/IeWUphNjmTIbx46hmJi6Jl9e29j3bgY1pEi9Wt7Mf99ZU9hCTuX4LfByMdjdym
WZrBVW+gHDzBT8YsB11+so1h+V/jZO0QRWZE8zZpxYFb3GO1QPtxUbsmFZyWnP7VKbwk83tnU61f
Q2zMIvxO5MbZaNcfbr2OWlHM7578JHQpBmA2uXUdGLvHBiMw8uWwgRNGXqZ0pyqo3LFQ9xjFAlud
DrtiE12SaiMozTgVuTq5M2PgNJjeSgxOcGpLaJ+Qzc6/60DkJhrLMADqZ5uaIwzb0XGg8ibqZkUk
RjY01KLiP/KcN8KFWle0PQ8li7apVvYatmP/mSAjmqg2YpPVJE+847cVy1JyU2kHrzs2jb9wAcdL
KK0VH5a3QlkmjpJWPNOjdTG223KQ9UqYJV+rwSvbM3WxjbGUz5eyy5oX9WxDOVg2mIANGsbpNlOo
dtZmox8Myy45/r5QGZd9zpcDMcXbRSN21BeMwrM9m1rAQ5MuoCt8kanMfnoK4AWHbdHuJ8hNQOBv
7JEI8wBBkuUoUfSOFVe0l72C4+psxX76f1ppwCbq93jCZuRG/YDGuyp0edNZxds/i7uexvKgunKu
hmdtYp9Iy3y09qoSHxVTcPeXlEqncCTOQ/bA7Xrb5HjzsFhYxyL9Rs9Uy54LRIYL5xmXy0n2D2fO
sCZ9ywEEEsUtwaq3XbVVtUzNc3bx/Clwy1bTvHapCQNqs5yeY+YrxEc9rGNkmOBdcVrUk2s7Q4Z0
5O1X4pM/s/sqVV1U8tSd3kOZyqyLVQdmzgn0WhOrHYfwn79/OWxyoVTrQXV/saMohC/PMgfj2Fbo
9HKhF9VPZrHxp8O7t6HHKPYUfOa1wYGrVNfyFnU3/a4vylGb7mOB3acD+zMkt7YqYgukLxbSMQnY
oxpMhTGCIgj1m93pGXX0hhWQParPecyazO1CJJuc07ZbcgS+ixMGmbWvPIccoSRM6hAGZZAY0xiY
COLmqxdB98vk8/2KFN/TnUDnt07mz1RoYESb0fPM3Iv2LvKZfrA358IdG1BXKu17yB7RHc6VgzXl
hYdwuZGYmw8clBVDl1+11HzOi833TZ9m0jlrVPd7EKKV9S9PIw4Jxu/N8ZMbwmghOrugDUjIaN3a
iHsg/QXV4QUFMr0OZpIqy/wHbhZVyrjtsdZgGjcQt/MceoU9zpmgFU7QQPN6qSnqTICbg9BJf4nl
KV0oqQQbQAZG6xDsHuF4X9u0FCVlmw2BwQrKeBvKGol5/hZ9DXfkb5Ml7VYUi99InLHezziXIBob
vtHpJ7c/nvNR6a/VIhWRRKTl4Q3xUR6Y9i7TGzPX9il1uhQSZM5kAmQTki2FMMZ8PtU2HYRJldUW
cjUrBGsZtp+ZhJDZ3pgB1tT394rirgwouibobGA8PbLVJ/l1l4+VB7npnpntJSP6N3hrx6080esX
ZKa9l5QeLqNisJ7uM4D8DULyjoQxiQIEYJqG6REDVrtDG1wy0D49PcoDakOrNT8x3hqyntiQkgAK
xNfN//dbRlNuCTveZD461+dwOL4y8tl1PEzSM27tJ1VxHzXB643N4K0yuoY5wPQCAn3kyY953p0L
48AKioV0k2dZZnUe9LUyuyWISzMQdt4uPwJD8cmyFDv92WfHq5UzoHekZmMBmV4yHCOkhFwZkb2C
VXJihOwJn3IokMIAIRlIBaLU8vcADpyobW6j7z+wNZitl5R360GFqH3yIHhmJnTBXBTxQAXbPC3X
xyS7gEniYQsAydGLgFH9MiFYyKANvfLHsc4fwQ5Ri9lesxYWhy03chHsV9lAoMfJrQGIJcW7CrKd
ZpdKWedY4quhLe94EPNjXMe/eeQLH3M5PiLh+kiclcKDcGIZJL3pqxAnabxtxQhwqj+jqC0EYhM3
2EoiEs+mm6yB98imutkjf0+fsrXWbf/8Hh7wH66aDdaBawnAfj4kgEmDiOP98E6us86JW7DBxb05
7nCn4nymnUVdIT51SRX/lGsMscNsK1aAFscH/vs5QrqLHw13rmWoNPc35ffiuEeXCFhTB18DIJ1r
7urzxyBQnTwtHBfYVCdMWBh0hgK2P1pZyYKDSHvvnXKFI6EbvI3d6T7rYbeiso0RQKi6HJKUihwj
CGTsCo8njqdwb62mKQopryWyJU/bux9bItqEpLt0+TAE3ZYGELTFoBVm5q+Op3SgXgc5kPK+dyx1
vXvgxxw5eBFNnpskuc7+lQWbBM14GZnR+UmOT4VhqmX0mx55OelUMapHbLHALqZLFGfB9rQLBcBh
tHLC8jbcPGxYNqTIbwLXm7Y76nNNtsyWC97O4m/0Vrp4lScEOEReDCdceKfIV3VEOXftDz6BS/1z
mOM0nuUk5bayEgGv5drMXmNl4LIF/X5fREJiIU7DQzsPdI9QvdhyIJabqae/yq1Z4rVyGvm8JJYb
ZjF03TETB8mfzPQhxZEPoNttpYloDYPgmzJGcUdcAYzwAodcUV0isNUmhAcfx2pwsG2vs0U+r4R4
y7UujUsZk6N6hXr+tW1g6uD0Ad3VENIgihKdNPcl963VvQkqhi2nZDYt2vgCSwCraUGeebte74d5
RtZ2Ofy+ZHSPHXHbnC/1FYYcoBqQNmhcDShVMGCd6CxlsGUMjYemSsRbluPxsmIGeSl34yOAFRSm
ioULf0747fekTbaJg1rXspPIRCGxAJJ2EsNUi4urckpuXM6DHTmvLbwY8E6QDV6UgglSk6ehAnR0
KnV2omUkDMC0JuJOEt2rHYTnLfVy6D79oF49zSNe2/ZNYn/f22xL/l3SB2X7lF0hALhlO9+hwwQH
GHtPR5IoMC3nclYNFq/l6iuealwdsFRctXyY6INRQYuiZGDgqcvRwyHfprmVn7aOH1K+CZt48pxv
LAKnVqOHMVHz3k8Butx3nIsRk7X6vEk9Kh8AzgdvxOEFgZTZjQhL0P/hgEYbBK3WB8aEK7acZE3Z
R9ohXqfSxM/TAnb7ZYGK/PaluhLxDkK0CqlCamNYybaw/pguYBocmhE2s63TWeO6q2lr4/57gWQk
F2ztb65/U/sgEkFRlEcIdPDVZ11ZrLgM/wktcHwMmUN17uGJzT0FLl2uy+W+MzEFrExE3GOvrAK+
2YINuUW9qATp7WMYOkTlyt7xT/YgWzJphvQc6Ju18G10EdZQZrel66KWGPxTQWEYCUY/yfgjlZYp
HDbumKPINLziXvUHs1/aiWMR4ClLCVJShP7yCHlYTmbLUSSsbj42VLrX+YxqbXnxSBN89oo4AUyO
fCy/BlIFiP43VvjIxgmBptWiFuOYTit3l25Kr24mzjBBEHE7sSL1Vei+KfRuN4e90b8MLz1UUWWj
Ykmq6qLtjTCbyTfkUGqM1fzPwYSzPaoLTeR4EyNBMfcX5hG7CiNVxfhYE+9OWfLoJxPO8wZREmKy
FKEgD+Cd0v50jAzubzauvDQT6+9OXbZQkiC7DLHB/Skc/JV8jeSTvwcNqXAZRyrU/WdBRQFnpOHO
d2oF/tdKHLDmVq3Y9wmrWGH1UZyibzYZ+1EgDupl8CzAe9RiZcx66R7RDXb/UUyl9ZjH8GPuCX1R
Rr05xpsydyIcI9vv8cn6F+fCtl278jirQw0SJAIm10/hq6NLu2Mj39lmW9bBh8Vkl9dS5H8Hy8uQ
L1Z/qanEOhx2LR4FqBZLy9+rcCAP4jGj6chLQnNBkFF5DbgNTCylzcdxM6OgxjyNt6poxLllhbMG
nl1f0MZD7rgMQpqPvppXmbTzAtDiTz772XPK0sd4PtcWvCCWfOERlu71unPf9PCRG4GPqggOLjj7
9nvdi79XLXGW9fpJxCqMBvUsI95oZ9ctzxEL4Fl6D3gJFFYT50VTtZqnNDhUfY9CpRhrY+KAi6sd
JdZniiGyqJ38U5FhXLXFLg7A6o2QKoRNbdDCuPYyvc02hlm7IvhpDK7i5ucdWv71+YCZoxetM1O/
fOrwKfZKhNQmWIE9xi34pQQR2eCC9kATRTNWFfIOHmroMJx4BcCxuNxmezVSd6r2irTFHTEGTUFh
F41Jmaab3WGbxcAHmmNDOt4qJvxLdGLf1YNtlTJVTZMFuDgfHE+voa+50I04c2gYHyXSKKs4/Ngd
hANAuPCi7PBOUNIu6alluYoHn7HvF/XlQbdtBWO/hM8uvp8Cp+ZPmyl6/mcmP7NnXNAFHXvZAlWU
eKHIMt/2YlxOAVPPtqnk1ILp+76jnYdpmoaCXkN0yZ2/0BjbX5xmrs4QNs0rFT7K997HsUuo2DAk
WQsLOu16N/dnx6XfSSAjyU5kUB/2ke4qMPe+PGR/S4+jfTpouWhRZX6wGy15j6iQXk9/LLZVU3ZM
0suBJ+OEeAKXwZZgw6zxcRyJKXHEHzXO20EDFbEd2Xz7pdVufY5WPffBatD0wkWLdNF4pFWpeYgf
voZ5lkd/1wVGNBrRbIHXhcrkBMRkGD7FvhcZDbV1Cg3qz7BslkOg6U4xqW8Kggjh3ek8WZEougrN
kj28LPDMLVjSCim6JhToxY1dEcVs5t1Er8S0l/gXXKuTEukQOo7g4sfMeZIz4oebALhBywAUjnjE
zrsGOlo3vqJ5PGHa00uelzoPXaM2maEFNN3h2jvWKh5WUe7GDrdL3LMNrxKhebtvkl0wbBvU2YfX
JWOcxt1gnWkJSneXrsTVe6/2DJYtshr5ARh9L3MUhA1eXSKBWXQQZSljMLsBFTYJo17OxAw2rVg/
I2j3sWEIbZDzTDAG3GfT4UEKeRrVqkSFlw+5RGxY/17vUswx0DCSxLrkC9TgvFbC7ukYl8jjo+Qd
iofvfZdz0h2+odn2JM4Fkyv9eFtpXW9cz8MFSPGFwJIzkP9qs4LLeagMcrIViOxLvK+fahYw+UcI
K0KDIwpcaVOpQstY5ZyUMpEH4cz1wh+g1EBqPpdQdJeOIqJqkn1T+sAUqmjrC5ACmuxlcEQOvK6N
JXcn/KZrF+bDRDujYBjFjDrCK/T1Ui5ehttUfqWCJyseV/QteajfYVoh6oC0d4xS+f00G2P5bXZc
l45mNSIpOzVfwQV1zhkxflbGph6W4YFc6KUklDOGjY2/toLymWkKr6NGkQUpwFVBaPgADsXM/oSR
Kld244yTgpLpQ9eqJyGbTFsaHSsoiQeppBvAcfqBtMfRjvs6BLmL07G0ktP5GmbaUfE4mJzAqVbP
Ssh9v7e9M9kHzG3p2HKXCHbz785OY/JvnLoTzmBB8KweDXjJOuKNJ7ba92Qhv4H+FOgdze9qgBH+
mXM9WYH1puBPczu46385av1Iz0e+Hw+a8xXHs90BrKP9RT73BC+8ohx5J1WaCSC8yg8LjyqeyiXw
DwMpWBJ7gxs1iVXHDlHMZcIAA+Q0AVisgoK/owIFUQ9mqOPL0izDT9eD0+cJ8RJy00lcQKWEpNNJ
MSdF3F3HN8nwx5TfdLDyQJ1aNvBVH9WK9AhC1JaBv6xspdJjLosX97QsPmSeECpScgiC6NqXjRoE
7MwcaUwmW9RihaCRajPiQnRWEStZkUe83I2chwKNcMEWoQPR/gdK6SzqchQIX3MyXDaolZ8vCWjY
JTjdGSt+594BenZ/vDD021YnoweDcjzvmrSyqzEFnbTQgKZoVQ68gzVGSHjA9a+v34VIPr0CK8hc
MVRi7YtMmqj0EIwMkzcNKLkj7MDXiFcNu1pKi/73Q4Gc4Q0g4EbDMBNAb5cGR/x0HuWmWfV3knuz
26GtW5Tn0jbUI+jtF1F5/pJTyeoUZlFCr34xeV5aYXVKxIaSO1aNl+ZYTWDdk34cdEe3cDdpu6x5
6+U2Z5sZvOqk6DOgLdqIe05A26xXgFSEBcHqbiqU3qHvLbujsenXlBoQ87JwWAeUiwM+SiBKC6vS
CyfT0esBr8IxwmZRLmxY1UA9aKgbQrNosFh5wa+ehig3wdptSdijAOstQ9BvqleFBaE9cLJuaO0t
dw44QRwUxmjIi+wnzLOpcuyio418U9qK8EttZ3OEqO5YHLCm5VYT6qgk1LH7Dww57B4x4Xsg7Kc0
9ecyulz8PNHSt4eaBGr30QcqOXZOdB6cRFZXlnl/3R2fA/BrWkDRBPCfArpy5fEBsmKDI2lOEW1a
VLTisVeO6IBkbCYZBMPmwMspvpVks5c7JbQZvqzKMqxLWNJS1bZSWObsQVOHv2x2hMcFDEt5czHE
M4f62obhX9R5EUtcUwvcmCuVPUefkFHWRqFeYKQZFtdIWeDsr9msxsJ5kfPyD36yAVdOtdYqhO+l
guMbq7VOuRjEfdwP4xolVzw7UUKmRVHZ+TIW6pxXLWzBR5suOtLEyofA+NBx5g8yoTiX61srYb1g
pC3SUIGidfL+AuXrp/yBSeVIdH7GhkNRTd+g5/Fkykd6hSdqxkksjDtHLZJ2FYV2/kzwVryKTBIe
KfZtB8u0I7Hs4bLGIXiaghCI7+jzlw0Y7ll53rqGuupkQmV3l9VKJlHRZtOGJkTTIthCYpO1Qfu8
vmyptJMR/2MDpvUlIXLDJBwEq4+ru9nOFnXNgLzguP0l7WKNYPyv7nQvA099H3xezw2F3brw1tkc
Hct1rEA6ir7mhvxVNkpmE1HFnmBW7UXVJEgqjKX5wrZbF5namjUw8Rv9Pav5Jtf1tSjYdURraQWF
4g2MbpIPDOHxspFKrTg2dzjMNIl9hywo7GTG35aUfj1uJou3sRWQtAausi5/3C+sly176cydwQh+
E8jJXFXcNJYrWXCFmYu3BWVCVxGf/lX90znQNt5XmtOPMydpGThY54YP+UW8zbEa+0Gigy98O9+A
ScaWw5oEdB5v6b8xdAb0zKy6jjgYxVo37oOcg/h/tWV6/it43rStBhMiodvc+jic0jQ2T+SjPw9+
Tcn3eiN3/rAU94y0Z6/zsMSSMmtDhDbvC4OdsDbhGPAJiIoUmXJvstdZWFHBToKkQvsULQRWDmfy
Gicb2qSV4Qhf8qT6TyMYIe7JlWEAkw0KwRfp+L/1VLMWLwldYr/FzZsat3OlX0vkJL/MOUhwSjF0
1GcuHTGgZtp9qd2FSTmwwG4df1FeSRfkZljRTdGToqV7lCe8cpZWd29qQ39ueqFGMMTbxP/MMfVB
K5iWbEfggVYFTNpqnHOCsud0PAKe1X5rj/xgnK8UGByJ2lgUTuzcvbdYn+oeDtpwyEhmv6+qd0ap
tHPtZP4aAZ3MeQDpH274t/pduKijobQXePsoHgREhX7OlyJ+7z+CGPOrZ7dHK9DSKBl7dWB1JzJL
GQLGjzn9lHG/uKFG6pd4rUVfDu0VBT35Y4KNxLjU/44eyqolcrtAlbB67zgngkFJTBZHioDSf9yB
nH+X1H06YnisdhsEkpMKg5aScLLyixJZbd3IGFs+OCRIGtXEADJFvqrjxMiEGgMuRoOiG/PV75Pv
UHil0Pcr7wr5Ec4UJwsMXyL60ycXe3S372ggMjTtfNShMcg5Frtiw3uXA8w1ywjYq3AJUwk139bz
Ls8qK+6idPQvLHu/jsP4CySF7stKpB9REK2pkz23/yok+8w0cFBHV1wf43e+wVSgo8mTB/sjB3RG
aKZdW4a/4zGmbl7XYlLkDYsEUu+/lK503TQsP1ow5g5aP3zZWvizHJvHRpfpwpMk2mTilcRFAZwL
GpCAwIMgtvBqq1atsIXtHsc7FsQLs9M+/tEq+iW66DFUhnwhJcWup6mFxnytO3WFx3TTpybYtJOE
GNHTaEZJ8pz00Qc140xmK1dLOZknDYUb2TA0V0XmJS3DuE+I5/uMEj1jYvpCkvB4gYMAJZ04leag
uzHD31t3qTOcS+gwDe6BCIURPMaqCEyqx9FNDZmOLLVJ+Ju1hUdM02uO5V8zWYtts79o0m0skRht
WbgG7aPR+vnG+/4LI7HZTc+RLyRHglql+ruLn18ko0aoHqUCAtwD2eSd2boACbhGl42EBQIKuw/3
RjmT4vdf+Rm3NsmnORsWjsYNhYScfK603TTaetjcLIJ0sCN1ikrQEL5vYyt5L0wi9PYb+70c3GoJ
rle/Q5orn01JXVwSj6M/6oN2iVPuzo/Zz1Qi1L4+jMpJvxaDruHLJWy+t1a8d9Y/xfaCxdV9gWHP
JgXT8MEFU4GSxgHGYR+RTiMQQK/uEoRk+J8e6CwTheWzsRbbRyBIHpuc5g9bOL+hlX414hfGTi5F
bogLUO62gfyh/EaxMj71LxAlOEOnHB7vmvH6Zga9S494PDbBTsX8b8nt83lsNd8S+xaBP2qaXGgF
SfFqZJbBSPfL5xpVPQc7D5wrLNnL9YKSipwElYadPaVSseouFGOGfgyjU54gTvUxMtNLoMQ3KIVC
ntMa6MdlpQg7WneYg2o6JuvHlCiBza5YzB3XDZBZPl7IXyQ42BX5zPzK3os4nhESwChEHc1oV8Ea
MidgmkBDs9lrupjAnL3sTDtmG18IUzqS0xrOYvrVAwudpgI4t1IFHmfLzSBCO6ZQluo3q/Gcph0d
OXPxotA5K2gWaViy/IUiNhYtYkzPuTo7k6cd7IA+qtpWkDk5/WEUlx4GH+wOt+kRmGrfe4xtz8uk
fjX9v4ydvrPLrSZrrPKI4R8lhp2cXfXDakjsjkvfE4jChAAiqnYb8VuL3dIhsjI5bBrGAPUAij9b
/Jna7bcQdXw52H2Vw35bzvptf1m7yDeqGPPi1j06aTDFQ4wkmBkBumPt+PBRfy/RAcviCgOh1E46
Ertg2dRXdmwAMMSZ3I2COor9uz65l9iGcljoZ32IJ58ORG91KAbqH2w2QKFbOLr3NiLQ8EHBZ6Xy
dGk1zSmS9Ltk00jfRRf5b9DIaLYpeH/4ZkE7HDqx6rBf+KSc5WbcSjrmBat7Hu+/+YzR0bGi2gcK
sOjXWpkJi9Le9g10DSIoAkUcDOEsqWp7VQSCqeFYVMTILL0tQ+uZQyT7fb1XdiHs8oFqsFOvDchs
g1CFp7f+ncAbjnSzIsCQugFrUv8VuAbKuuJSR6A5XYCGJV3CwIestisaqcgrXm5nAX3QBSafSAHw
xb+hnbvlBd5SNDjKh+MbMA0dJcpYU5y6UD9wVTbNFZHL7TNen33tjMwYHbHBwBD1A6YJRl+9nYjP
aYfB1/gV0nlChs/qwHYdaLr0++fV9b56VdpyVDEdm5TbW4FwUOA4km+GOKJUMi4ZNX6tLBSHM3nx
zQvkU7lb3t3yLVmS5hYyS6S61LUVHAhr9stZLL0Mrovxhx6UTZcsNAHVXWTJ3dMe+8wEgZFe0pHa
Mw9ZyUvwW2mnUuqfOpGXjNin/1lHnAJoqoBNOazJHXaYSJAf3PDK2NNYuF4J3ROG40eVckIlFD6f
18KdV2SZCmhD8B0QDLFduVBEaF8nW5ph4Vrc44XMKusEznpGz73ZYSeddlOhvthTPLSEfNbs/3Jh
iySHuVDARrCifaUm0NneM27XH2Z9wQm9pVcYLYCclLSIlZIKcGnbR62D4xN54mvWacmmnZ6D7WiL
cZYR8moBY/ZMTmG46Fnl6yU9jcyFu20DQHwIBRRbcbS+wqKjN9p1PAK1N27Cz5VH/50OgOn4fdTW
o7OXlThPDMEH6E/cEqfS0ED/IyMquzs3KkIv1f7ZsBduNIXe37n0+FqWAlem+y+OYNbAAz/ABGRC
UJHz6rUAaWP3S4zglYYSZDpmW4sYDpo7eBc2J3cIVxpdRJpTKBEWfTl7CcmLsyfPTE6USWNhi3CK
fu6572W2Edo473VVfI44uIc3qER1uYQdSfetD4iXXB/InoP12+XGkVvqcDKsu+ZXjE863AyLOuyE
3Y8UGHO54hJAPz9WNZ4b0SbucHAiWvMudq29VQWgu2hy42R+SlQz+MgwcEld47AcD7/WxJIzBlMz
MUCOUEvkNpiJ1DI/6XqDeXVUMtqQWTxdJYHyWWKmkfrUzcCoFPYesmiXPVzcgrfch/paI7EABHlV
OqMmInY3hxq0jLy6ZpRGC5DatFWo0375rf+p4iigXVCaM7jLD80qPi69lHPC8oU/pNxnCABOtVtZ
1JbE2TA2g3Lmaalkf60kQzEiGwU/TvuP/219BchMvA99KT6Z4KQWg/BeG1TgCk0zXbdKEfoFz/e9
uAuSFwplZuLVmuvA1I4ly6O2FokLexJuyUhOvPLH8XrYPzKIMWEGVa9ZnqUJcpCnRDIdGeOYZAbZ
5cgs+W4ZfvC7dY830Y6vBaDbLXHuFNbxEB/AKhfgMjvLjdvLIQ4B73OHv5VwHOo8GABNpg2gV72m
OtjDbresFMejOB3lhp8s2upl9emMgWS4V4Fu1QZpQEU7D/W9MRiNtG5H9Uo1ygDpvBom8x1cW+i/
UA55JLP7BJY0ipPmDBw7RJt1s6AGx9lDLNAZ4MBglruAIPgPbQpcvuJmp7YseqGl5yFTdh3xI0yd
D4TPXd5xaIGKtGtPbhkZIzEdr4qe2rBaJY9gJdpGuVZMhMj/2jnuhWMSgeosAJcOcpUuC9WB6PRp
h/+taDuk9+TiHTtAu5/9iDs9G1QTDa3JvVo0Ylrf0+kYpPIcR5QkyD1ByKClIIGjSM0BZISt0LZl
rSf3FDRGd0BNDeKpxNL1bqQiVqkHjiF7SIDnz6WsuohHQgK0F5I0BA4ZEHnVAgTOAmp70wBF4VJN
Gr1WWzSyU/epdY/oC6qkSa3PCS/q/ZSYbYw+GtcGiyPfugbdJgpBQ5r/gt6gkm3EeRQiYvtBRvXe
J5RRXJK4QLyDwTJ9jhwXrcvhNTBhrUQc8W+ShYIIDiiKNn1A7rTOL9CeFPXTitMuXGdiBdEb2wsH
ab1+AATCnH+/Ix22hmMBX7itFNDVOgMYCi1Gofn7KhW/pxX/1jGOqcw347VftLafTHsTp+RP9q/x
hldlmx7dRw1Rgdb0BOZblXoOXG3ypHsDPRsBIhMJiO15SgFMfatYu4sFYb9XjTGog9P0yl0l7D1p
febZqXGyD/6p6CCriRdqwQQ8J83ff5Pz4hzv/3DOktNqh1X+SjEv8LEMYCdctWX2AbtYgxLBdsFF
b58Av0Q68cLLJ0nJ4ZPqVpLYLDYinjKGuf+Gw/stwhQbWF9CU5xlFSs0kSghJvc0kYDz4Z8adZbR
rhRq/kNyEUObI6wprbI4E8uU1QZd7pp8AoIqkYXkDROx3GhJnvL7OxIN2QHBDbWlGvhliJBaM6C6
HmIVmfmqunu41tgwSTJV7aPKekWDdcKsyVqPyTUNo8JzA+sAUQLakEDhC5V1eE1ZxpZ5f6492CS4
C3PqXNiJM66cilyxyFpJFP9xff+zLXK+0VH1e6AI19pqsuTfdcIFhSEz7pxUEPzDv4Hnn+O1fHkV
5za6vSXoRqd5sp+RZqTRut141uxFaI62QKz33aKll+L7nwIefp6vcp02xw3rhURmlAZPLm93npH4
wJg48CYXCO2wORmr0zOtVehSlM0hOhgI+G1R6Jy2KSJ5550sI1BMt8tWuipBuNgvhfgf28EX7HP7
NEaegDLsbmMH9bVSxnzFhKSPsH7s2EfVjNk6nIDQrpiOKMYHn3wOJ9DZw3lzqcvYxYpEqyvYml33
zdTtVbmUAxKqQPn+uAWZQuvpjfj33Wel4XLPU/EMAmJE7Rd6i5utlpsF4jAAQUNVSN3hamXFO0J1
uyVmN8RQ8y6DnLbrIC+RnVSJ+FYbj5fV6MohYWue3OM1l9mE8LxB3zOaNWlMwC5srXSFL/7UjxLG
aKCIgVGebBlgpnzw5NuXOVvFa0ekbjrTKFjRA839DNYJgz5aEfaYtBeiCt+Gna6fyYXzUmxSVg6P
2wTSUHcTsiz0KpVQH/LRjYFbg606fTfFal3siXYhUoCbdXDjIwFeZXroGeaVLCAr3aoyJfWDq2ex
OemsT2fflOarfQcLUJQ4HIPz+9QhU+rVK5Exv5HoPh7u9Q2ZzJU1u/N58lHxiyL9UyYW/F2LQOu9
jj7LSNU6UyjUr9afAIsy8sK6lIa/FUYbmQzmgYnqtwGoRSxGDxSzSYac+CuQEQG8kOSjrALbE7Jy
bm7fOlpbEJM3d8Ib2fNIo4gzMELXvtKQNSe+Rmi6BQwJCx5k35WO0cKFl5zEJY0wte4KlHZ6iuGk
ddl23VL4R2sGBi5AyimMm3cJNyV6YElfpsapO6/qV01zCxbsCZYqQcZqLfNWKWSyHpwohNyLLetb
ysMcCowEYVIEwsC+vmuboGMNTav3FAQlCiyN2fdLTDjVa2AEZZe3MXtrKyj1lIB0Okz/0lkAL28V
p4a3xWAgG9tAEY2VNjsXyehnwhtuiwaEvwGHPYNBNUo4zG0lV14gSiQwP+H+ZNNABpbFTXjqyiUS
rhT6lCg6p46O3xoI22/3SA5O7cawdBECUowmqGAHvuCt+Ce4rkulDb7axX0gmNd417vuqSpQKE5S
5uFKb+LsQQ7VEEDbiHtl3jBjZBKinWer9Dx9YigGzu9QJUNeK85pwyMrZohzgXWrJwLoAfuKjkh2
5uhg14jvjxEuwlHEAHCiNJ/S5yiI70L9vcxsihbku8b1fZDvPpS9VhJGxHd+soxbD8C7G8gExu4j
xZkvj9ckSHzW0GhOoF0coinAi/5RG/czE0xwmFuEJ7WzB/z28xKs4qy+CS3PfXO1fDUNHDyOVW8T
Dn/ztiKMsZ2myVioXHIOuAnx64wnIMj5Dbm/d6/azkhT1klnVdSUAnFP4oFbfG4H+VLRY5Sko5jX
1wLBy5h5i2fa1qTQxYJZ84if+6lkCwDb/u0lApJa9zRMUowugsU3CdCJdLFkiov6Gn2cw4bAH2H7
nDp8JIIg3irON7kf29iJ3/uYd8bNXZGj8SC4pr3xJFHIjVN2dY6kSWw8/QO/+vJ0tMCW1fOoP5ap
WiB8k38TLrLVIrcbBk6jrQrWCgA2M03hp8MneEEPAH9OMg7StcfOiqxQs2ak8RfdC36gfPhLlg95
+kb45sVA4JWPioot7INKMmeV4P3K3DgelU0gVwzXAtwrII5qRtqFCxQ0NPXhrg/hV04R7sdqlduV
qDrT/5SLz6dqLhqDVnSHVZENYv7izlR/d1aR+gZ6tlPm6X3dt71LZobYCzoF2luoFD+x6zd8ElsB
gBG55ODUFiskDil9CcaKxChbL8eQaNKInJM/SPYGJQIuD198Ldif22iDWJQrmln32y4AQlKsTyqT
hKhYgfha1sM6Oe1djtRusntRT39K5l8xRMdte4iPHa2ML2RxXgW4druL2mZaIeYsc+7pl6to7kJU
oyj6MvNXXwnoo+uxbGOxjvTNovC9Urhh7403xerSarMC/ZPoikMk84dk2B7rP7yvhz4jhJGnGALm
8+OvwcmxXIau4oUKb4C9ljgFwnSkGQFt9MLhDBNR50NwbtbTYDC66ezN6lZkdyiaAWprg86HxImE
cGgkMMJ7YE5Q2YV8d1+ddolvaauOuQNdkF5DslkEGE/1Kva/6bAq5a/DGf+AdVWJXiciQA/BBK73
8jsEO0y06c2oj0RhVxEnpVYx5HSpLs5UW9v+B8sC5hRHUqkoTOSJi3n1yKLGwWQpMuqoOB3k1tJf
/FsxR6f1p/4cBYmJyMdgVGWCx8Bz3Ngs815qkPIVjB5p+f/J7eScHrbNQvK8bEgoT4BWikpF4pIK
MeGmeIBdKck4xie0A43ZLhXRxtqbTOm8ATYDNIdFGGjsLgiGuw6kMIEwKFVGDUqPlFSQ3yvhP8el
t0zYeZ031M1H9hI6NmtoIWvrG8earsjeS/O8sI25HiayZ4Ij9Uop/DAg9pNy7L2cXYCLzpLdn8+o
gVrBRa4UEcHwnqiaQalFx73nxCn5Mhm3sC9+Bt4NsghBLjzCWqcLSpD0DTq+83gKJamY9VCBCJIi
YifHt3IiT8Z+t3zSO6WYCJnGgK4fwQfj5fdILbtKJ4qYyODOnUqpQ3la9ZzuUnyiqK9CUR6vLcCy
lEHOCHVaLQ1elUr8Od9aPEdtrV+yeaDsDIokiusGT3dq1iBfuB1hjnlWqEDvM8y8ZKu9MR0D8hxr
iJpG+WdMSx4QYR4bv4XlARSabrm9N7NRh3aT+cYYclaB0sPq2hGHIz4HWDhN06J/AvJc/+5AkTpC
b2L85ZUAEYh+RZulCCzQqrDLf9bPS9KcxfZT6F/+trIpzf2kJEKu3RhYz8OzE7hK2a0Z06fYVbVT
n0ofVHPQhWZm9/bvICybZBBvJudy5ZJ3aFeO94/u2RF2STknpdM3LiDrVtpLfnSMjasfKOwC8n3y
gUnaRxQnyWSbib2FyEuHK2jg5Z/IVsQzTHMxyZ8puJ9KtV3Xz16lZBYCPyj3gfoTPiq/iM4GaQBW
PF+lznO0TS6sJ2A44Tq25VnO7bj4Qe1BMq7uYYzBhOsjJbwimyPSLtZLb67ejpz73KdZ8rJYMnH9
YrynzyDut8ZQwegp8H26xcC6CvhTdotna8vq0CnAc/ArJGQ9BAk3uDqPZ16pskByzhQZf4jm/0o8
GUN4o0gofq7BnnN0hwvnNgDTbtrh6S+sIDDvh19uI5pGdqvcYNGMiwedclppSYVaFmAj/w7N95vY
wiP8eKIKwpK/nSmahm+HPkZZzEob6+TCF7U7n8ZSwgP8nE57DgHWka6f7YgByq5sVYtGOKpZijft
0YAy6IQdwzWn6XudLDPKOJpZnnsZLnD3SnvMpIt8uVOZOL9mYNmF7ZDmkt5O9txGdELHkOgIB6az
TjLxy0ytJbCejkJDoJ4qcV9/7+GLlQs1uPYJ7N3umNpINqvoLf1D/hy3epfTh2dizclpm4oYGXYu
38IM6vWbQPWZhM3fZIOvIMTgrcaE94NXkBqPl7OM81TCDj8R52tG6TRNR0WMk0KlToJHe6Tk7bdN
9zE3J4a8tbDdiLBFx6DSN0zSUf/jZRth8fop25NV6BLU/QEiRICMioMd6I686fBEFiUv68xgvyPZ
zpnu83uQjb7ysFDUvUo17bLf8AyPVH5E7keaXLgIzvtoJEuV90h3Wlmh+CJ0HvQ81l+2kne1eCP9
m7hI3ekmOSsZFL7gn8fehx1eNGhtMGaSbnw61pwe/LXPIEpqpgOVCrqwyyjwz0JnymuxXga9iMqU
2UXubr+7ToHY3mCyDtRVbO07ia0AJS3IfdW+p5xqfUmg4RvUVmVCTwq76bu9PKr01pDxZyp2r9rh
3d45XXFqlMIVVWEr0k5Jl3D3sI0hs9BlXSF7DoAjLox8jrAtMQO3rRE9MFSPMnUmb5VjLj2Nl0th
1XdPHGkOTT/U+qvUAB5Ye6prUJiS46+8Dukexwwojdsp7tE/9ZI/g7ErJDGwQAvbel5PJzuYx/28
fo3R/VzCtCVNY5oKIJZ+x5c9tqwMEwyHWDTc1IoyAeTxQX16UFM57KwJMNXDKydRAOMQfVaCvzun
GBBGxrAN18gAi2igj1PxScSlWe5W3VpSa0d1rO9CLOt3WKNTIwPV99z7J5nMOPQOU/0E3xXqSr7G
RqSCdYeLy8KfjYscZYSG0QMK5xNwwq0c472zS/xaudWcc5nSEkhWahX1kK8zqjO553D0ImibpUKi
quPGv6UHi1dYpCqE9xDB6jDnMwu9zE1gTcdKCfvpZoBDfHlxKbEVlMEtTfQ1icSXLqWYX6fnYNnS
pgliqarPFGRoBeMtrC0w8VlDVqdKAbZKvag/9EJ1bn0ukWF7wNzd55ssW7vIWvwyUHW8Trombbsm
XIi6jWJLLPCt3twqxhnUvAzvrPOLrRh91qnp5UMN3t+nWdQX6PazzospLjpu6UK6f/TbXzBdTZgR
z2Och8rREUZK3vKjkv1sYIvE25Tv2cFwEKCKopCq1mlRRz/JYAXzi5Lqaedd7zsOSUdbb6L1k/SU
3bC4G+cEv8hGndKijNpBij8b/fCMaUteJdacGWj0U5r9Ep9PjwxKL+/h6hPzuHEymZwGWNDcI7jI
v4ylKgHPB27VEn/Ycrp/jXJgdZ0tn2bETMhZohmRYkYE3j0L1VM1IDvQSdjizoChhSAzabJte+Qp
KcYzbTONIvXgArHMPkhGvSLJvcf86oxcc3jHqYScbTM3YFrJVwsU2nD1q+9yAmu997hzAZFUu/9N
qJFZs9lHxW6QQ3GvISQ1IjydCeAaGxr+N8MMSCUdLxVxR1x8LROIpDyWi4HQe5eC4Y3KCaFTW15A
2Q+9dlVwM0jmDGGktL/sXQo3H18jNoId/y9nlm6I8nqtPPLTXevWmTObMcMYx6jsw1gnjPK/dxWq
SPBf2lAwo8y4nuaopeN7Jl+dRe+zDf3nkS3qXK0oEm6CSx6X3lh0U2bDB5Hm9FINmD5wwqHM5pA2
6I06F1pJom/Z5oWwKn71VFQQXH5UcUj1JAwdkMnlwalb7bNHttm51IIpKC+cmuT9FU1Ts1cCa3S+
e+LbjxMzrHv+XCAVgtcH5JGhzJMSKWx72MANSOmDW0ej1JZr29/rXlyc+QqtlGjqxUtFxkfpjPUd
N+qRikRvo0Ug5wuMvD2uz1nu1T7RKvYxSyKW3w/i5l658yEVsDWqZPKtcgh2MV7Xy/MSouz6qSER
nZxYUeIvlNjq5FwDUq75vaSvRklmU8K171QOfXC+dJWBd5o7WEjanG7dx7gk9q4SAuS9dxgN8b0d
QyATt4NQgmKEQXAGunnDPzdH3Wh5MWWa/ZML9OP2PYBw4o03V1VLzb45/XVdoR22NQ1ZV6xaATbH
C+7RV5z4CL+nmK+UJIHOq6LpXn6w9Rfc0vtnTHOggc6RymRLMhk9IU0Hp46KjzGXPssy53ZdY5mR
gny9D8NDExJmxa59RYUfPUsdtYNZmWOsGVM+it4/QPqqwwncadzfzXF8Iyg5ZkA0ttBYEJzS9VFt
qlKc2XaUs722IlAkJiFiFUwEtWrs5kznguJZN3+s51KBv4dkqCAxGrZp/5qD5holK6uqFWyH1KWV
mxyvhZOF/Bcf9b7u30vtilNYtpRpgbo+0i1xHuppOcbOHXBMrRzLwBtp1RBaii6OmSQ3LFNcIJsk
X/WVgsICRyXuCtvzez14kPHMZA4i/b3v9w+YodOYVkPnu4EXdMR/ZvN57pxFA28eM+bBgEnNjKAC
nGCFpE/Xc4xb5KBcWFVCTwlBRIQ7G+XZMgQUB7fxIJQ5gbmvR2jEEFA4B0DXLZsJgXg2KwhE1qUr
9cdgdEUTPnn1A29wVq0Nj+K6RRf4d/bvLSPbSyPn00GbhWj2wodKJql7HgKu/hbEHYYMag6HX+PL
Ym0Bus6+Dj/n93SIzl/D+YSzBdaO6T422aGHXVqID6ie9BLUeto5tSZJZl5xVy3GGdjh7ysgRVcF
viAahsbV+8mLjpbqqBpeEXRoFf/KPBbJtKm9voNgmfeT+FUnqqBpxXnBR4oed0jlEyRhYcX3gqCs
Y6AIvtsB9kkygxsLBMtruOJNh0oFZzngN3VOcnkECyHmWOPkZg/K0GuZ/cKtMlOctdgpEB6Px3JA
FeUzzl6dTo/5/lHHgNLwp9U3HUOtGBcdKmQl0ORR2LAKorQT6ypj4mpUYrzBGdfNhvL6phlcmx23
kxTaALoeVIVA0GHDLNmxm5MwaHrgNDSCI2hHOQoxqxDQS51fweJo9sI15YwWhYjp1vNgVSIKg6wO
6zv03sb9/qWsqm/VvDCVcDfdKbPzGh4X3kA37uonbalVv3hwcg7kRP9iEadh9KiInNSqLJZsL6mO
S42zBTd7AHqkmWRda58uOLeR5e/0Rm9uksyGxBwOJ1J3Moi5Lu/5F4Jxd7+s/35VHsJDjXMFSuH+
JvvVMCbU9KmPqvHxGLhmp7A6SGNwIjkpV9E+vaMAE7GlgYRx+d9SasTO6Ura6bHWoxJS5FZxsclN
8+ZrhA5bYmLhLZz/hpVVJWdrUVcv2S/jSboeu8BYlzVKsX3Dz6zzZdKoKDJU5Zq8ICbkoCrD6+79
vsLPVWw8jx+tqRQyWrYwrbKlHflp2gwOTD/2u8uY1hszO1OFdv5JfithWIOnWY9hr0XHnWnUU3AX
7bNEYI64//YYgyrPEfALR+mKdgkduLTUMBRcSHRPkbxVeTujnINRNeAgitAFZyZNhOdiYFuKykMH
W13kzDhe5XmiuQzFdK7Wd0uI34s00aPPqg5DY6MlRrhjg+sDpJZqiVp6TCS+FYW/GnowN4QI7osa
G+0kEAvRe2GGxxeqF6u9M+0AI9tdAsm52nBn6yK8y0ErVZ0oinTbAiSSZmguSibWjSOufyO+57Fb
xqqXVvHPuyRam4gyeD09dHYJ9Pg2JfOcMYJ9yGLiZlB5kSvhoECHl55w5gWLHvKJl2UiuREm43ie
StQ/T4byOII6g36Vg0o/7Ctm37HXN5Zzg0meCKhwhyEE0BMYpT0o6CsZOYZlU5PBbMgqhgxZcpZ7
1FQHXA15t0Q4c5T0Qv1jLkTGCmre9dF1gvRa/c5s59mM29YPDLF2lAf84vHlOpm7q1+CgfIbYx0B
rglsYtYp+iD/zPpGw59Lta0NUB+R4Aa4w0Wt/4dUww1LwE89F8Jpa5Ic183S0ysby4o5uwSOM9Qj
P6asSuRb+9V6Y5/pbVPovF+AKztzxqm6rzvUoM+zlrIppWcK4blGV/sD/41WrI9Rz0x1gAXRgJy3
JcgUTeDMDLfLlIvChiPDTckRDcB5o3mULmxj4IGonxs313quNZshvY5Xx51FqHHpHZaa68I2ZkM8
znW8v+0QEtRytf++umd+nzJk479eeis9yRtOUL2COpUCwh+I9RvWNM5PTWOiihpIQ17ptFaPny+B
J0xzWfrGtixqLZGOTOHg3QhAapQPTyKYdjx2XZ1xvIGDBimKqjiKvV1MnsLLwgRS+7LzzHed4CKc
k+YxXSnh7gOYnil04cO8E+2BtKNGLajXPeuyDMKWDKjSkj6iQMbUpCTo8oXNpZ1wO8tfGz3hQXRp
ozGBhuXuMH7OKyZmBQ74DrdDCCgTuCCx1aotETnHXBfn5QkGoqWvBlzYbmxvXWpqEnVpGWPhC+9T
s2KxXyNnB4NQdEWy4d1s62VXj2QodGToWQllOWyEDxPvk40g9b6LvCFJrxrCbodAFCfiuIF87DyR
OH2F9xlTAGf7KkME0r1BIJyYZe0haDoXjtiiVuhrF2OiRUdlVwbxOLVRM6S8681XNS7Iy35aEX+d
vG4W8y996YlGeWZnx7TMEWL25zWqnCjAXTDjCtSw9tCv8goL+cN2n2opcV2wVtqO6YWv1LbAUUhL
wKs2S2vN0ZhPcMFpPmCepHuaqsKY5KnOjSr0PS8HbfTw/xymiAkgA9iDm9T/WfoxhLgZ2p8q1xf3
OUVyoHy1RqZ3fLUwO7iHUAqhK1iPlaVIsy/hfKc4vKjI1QT0wmxAlBpPeysHkMwACtQOxdSp0T4y
bWOY+IvCiiWYzIMPwUB4onggHbhCYmvztC9N1UOnnK0B0QbH8a1HwrZKnE8RAPk/Zhh+COis4lgE
mssEd0L97dmYx4OCpgmazb66C4Mp3aBowngLiR1x/8EJiBEPVnCdeQ1pa+c3kyCYjq1M8obuv4Ut
UMcVQcWNUeFgXUmIAw4o6BU9p3+ssdDh1VkPd9Kgfu66tRJ/lsLWqTIuXs6Q3/64szj/zV5IIhJr
iO4d2AWe5RB0lBOePBtnL793m2vnakAQC2dDzlDJhK3vUEQEz5XnRZHFRw101QZhOKyk3ejEJLYJ
xf5s1pRO3W3Dd5sk/otfR37xFySBk3JrXSWzfIyY4MADHH5ZkPPXpfqv5FUym2M8ovSjl+RzF4dX
h2jCGcQrLtAja8l79IZ6Cq6l6m67+zReoKBMQSu/7EvUS8PW1yhEJz9JXrGNXROrDXuh4/ie80dN
NfRjVtILV1MhqmIzXvW805zIDZW3r/ijOsPWlUHl4rHayoS/o0uA2jSEv8eBHeD+2fgQXp5pIXQI
GTAWvzmgV9E94y/LzGKoyhf7ASzhqKwREKoiLTEtrMQ/3spKjjh74N1CrdAWeh5U91rBVL5zOK6F
BwFb0h7RKDaIk9dgNu+QK6n+ngkbo+QRMtvQLu2HcComIMD/ppN2o7kugn277kC5prqKXAxakIfO
LZ8XRztgtw521LA67vX5Gf52iw09Sy+q3csksQiaqxGHJ3e/r1dy/+WsKSEa/6Vda8mbn3iqUflj
/YG22fuu0kLmLx8F8wW6U+vwg0yLQ72SVRoc43NwBYSmMbAcj0BIiWld0ooPDcGlkqOcJNQtQOVP
RZXOLRm1kw5Wn/O6iYaEQAH4YLCWwWp3IwER2F3MgGT1xyO4bGYtArBOSWEZpD2JNmj9CFIn+Bqd
bpQywSMhoigfWn0oY/tukORa8mA0cXj0PJaO8bLAAbAdFd8l08FXbT1mLBG9tz/DYThF/wGBluYe
sCpwSmqAyPxHCfTYogT/nLBb5SlmWO+bZlNMotWCwIHDRpfKI+mZkPqHiQMO2yVxCRy/VDAReiUS
lC1NNGMLhD0Rki9fqI19LU+ugL+KYM6DT7BKMO6ZhKqkZZJFpxUAKNr3Btecg4UxgabE6mT1vxhC
iHSrBAb+gbeNsENSf+sO9FQ4q7CDpa4OqbTjUF8PxLPTthLfjfs+BtiI7WbtE3ed0VS9wzOQ0NAG
HDYvlnn6lchr9OqW74zyRDQ12xVBo41uWbZYNMeYdq6QEqmOvQfal81gCLVqoFFVV4DAyQm65Jx0
v8uvF/jWXMZxHqsA3fsX5X4wlQd4HWpMxbJXIWKaHIW4w3pWZysf6nsZXh50n/CcTUlHphJyWE0v
SG5BMo5cE8IV9UNBx3i+Wp/Pp5gV3NysPfqFdtfGbDW2jUAjmf1qv3LuO4/lgelsl7FR5MV9MPqH
iKVVgBEHBMlIexogNlYZagk2f5w/zp7wA/v7N6KXSZ4SgBNtKWDSOicv6dSuli0xgUxpPFgTB3U4
F1fBXaXkcNUCyx7bX/kH3cuFIVgx5ZM6lbQCzxgrsMNTIIC1EKeeMCr7s3/1Q0kKEyV7XGL8s8XV
L/oPa8z0Cx4qSys7L0GzcwerREYBltL9309wIZpSfiG9wvqv6/xHkXtfhB9KZxsmvTxrT4bX7hKU
2LBqOWepj9Wx7+m12mS92Vwu2xwXCjahuqxCTG7h//7XAIrGFv8tATCD0fHXzDpocTUGUXq6xuxq
CZO225ApN0sQH0m9OvvpahadtnCp85WHEB8MGWKnnFUKgsh9BZYFFwBmD4Zjg3yn93/ih7IruWFc
37cFOtnqOXpnSmXaE2XR9euxV+PBqc99yrwpfo2ifOLEcqhBW24upRzkGlopLn1fssviW48IZovc
wN+EepuLbwlnI9GN2UZJv1r6+daS63Q1E9dxhn098MdaUYnJePkBa4TRt0s9Vafml+8oDXIqtkB9
0cejULu6qDSQ9LibbWqgLd5owTGmAx/jjow/UhtXWOy9Jx//WQ5rpYOG/Mw6W24ZYn0LL7SRJ2TB
b1vwYzLZrhIC0D9LjxsNLanUCzkgYrBQGC8n2wkayZkkqMk+kZ9k9T7mGmZKGmiMIaB1QAnkGPax
pCggjQFFFTzK0bHx7rG44bV+otnzOMCIABXnc74ToIOpCBMeChyFw3f6qwkTsuFIoE9vkuz/gkOF
UiqpCBk2Uytq6EwnH6ToZx5Y2/sYuUOTyZkF9MKb7qE1cutyFnwvIhv9JhIDKXRbI2Fk+bA8YW0C
+qvFjZfA5HA9bFTPBlHixwl2GAjy9VgC2amafXCSy3ciic1ZFAMxruYMe/wFUM5Z9BsXBCvo2crY
iC4IVQp6aoic11UmG+UBc38NTZxmC9i73HSZuf4UOxTnJ9nNgyMjkGLtd9gfbnieDhrWxzngAv3x
VbcxdXEc2TFPJ4qAU1VJUJ/6MOKrSUHi3oGSSnWnGFpLL4Mr4g7bRENxebCUGGIyR1AOL1jUBnqL
719XK6RQmTYcCROHtIeRtqjdUZo0sLyea7wtx02WnlrDNLqJEtWUB60wmb6o9/y480Ee6AIgQ7TR
KQQIjd55jYg0rhYiInOguluWc2dcMUqz2PKX0lXIX1KSfINNmyB0MiQeUGGrSiI7B+MpJY/ZGOAg
4z/K7NEgq8eFmPqFp4i6zT4nWqOylNg7M7Y+3Gkhsng17+J6QE+wWY/g61rUmegpMyPjqb2S+czB
p0GJjsUwmDUgKYioP1QTSgJ2asA1NO7JUoxQiVkuY8+IY/i3qZZCxBpABKMRQajVIzCIm2suz32A
L3QKREuSJ25vWkmq2JTm+4OnnBdMLZwY/tZf14FtH9MCMQJrptYYXdDuPlHyoIFAMYCyX1Zyy8Bv
PrAmymeUjD6sHOl62yKczsrQ+DDUPFY/HCqCICPqGFTAoL1CwXI9P3TAkB2g2heSc4dxCRPWKyt6
kPWdp+RxkEAMmNd7oklsSZ13/AvPCsAxWBOGh90NwEuTmx3zQRqdQdU9wiliMttWjiGBwV72Znla
WQDcX3jFIEOfT+iiTDa0YtnhYSrZmoOlabA0SvU/5QTGo1Nd5kLshVV67G6I75FAl2p9bIlMHogH
UOotPWNFujOg8BOzdbpkyA0vm7Url1YdbzeV1eRuGCZ9rJM+vNfRjsd5OsfISV79hIXpcPto5xBv
b4uxk7PpHxKhwRX+tEcM+k51NuXbmDM3x134p/kBmu/liRUSL1agX0lUFQpqejjHdJKRcd8xXeE6
EK6SGMJVD+67qKsaX9dBXrgNlBp0Oeg6V59MZPJzqNRS7PYa5RBEzDW46cjefGUalw5+nY7xvKXn
w8dL+Csjz2UD+qlm32ef7uGvY404yLJxBrxM+79vXGfEwX7tn/SQWb1omxPZ42PPn0aIdRFAWOQy
m0f4jqRggfV04j5C+bCCD/GICAzKLHrzC81Q2RsU7HxUljwrzGGC917xb6EaAgOPIGhejZ+lgJzZ
CL7IKxF1/RlaIFCGv4H1vPzdTy+N3iflWAMwOCpy5RqGgRBQW/oeIFToPwqbV3fI9g8n+4DpLvRp
u8/G71LWrDzWlj1KnUyuQNI/E+gKqkq5R5GBbbOaatoF8Nj0Kf43JXuWJFvVt/JOyMARbMsLelaR
maeZFY7ZV9X1aj0fy69x7jJeVMXN/8kLxK/rUVP29eWQxs656CTn7+e5tYffnqTIkNCYmLDhZETd
kkM7FyVRc0MVE7whL4hF/yUGP3ttTQHJdVwT/y5q1CSFbE6eyNKFj+P/wt6U/wIh6PLM7r1BEHgo
TmQczjYUM1dxUcfzfSyuIJMxoyED2eirM/0gJ7yYiapg35kDMrvh55mXug/w25o6CCrmUGQo2vki
B8lkuPsBISQpi1wjZdf56VQDz8YC6TL1TMBMEl4b36cAvsFFL/jFCD1EtyB+8ritbnCeoDCoH9lQ
fpeeq8LOMjrhTTMIvI9epDHyJQcwXl9KQoww6jMj/EoY55RdSGhgMKS5MXyUkGR3f1FTE53KYZNd
7Vh1BNR9C6Mw4eo7RxsmwbB2rK+og5hW5NdOp46+xYs5KnGgOsNJ6dBFNu0kMdevPKuGloR7kBFa
s9mFnvAWGx8Fo9zjO2uehVXOMqF0J0dFh07Seyvt+AZx+6oo1CAuftNQD10aXDZQsCKZENAihiM1
/m6TpyHS50f/BitJJ/C0NO9aSVIWr2CepnZCntEsC97B6jk5TQpgpF3SGaXg+RMkd5eIWMTvtJYG
CX9YncGKywCM+0tO3+GSBy0O0kznjpGxFcmx9yJE5pyYcDu9bVhRHtqg7YmCx0R2vCTpu3oE/R58
ZjFADrehGqY/ZFfumFWgSngGFI5h4zCGpWHLBMb2GsJRUfMgnUdkkY9RrrX4+9msvOlW1iJe3NMK
h5sBL44oNuA37kJKfjB2lm8sl57D5FYttmlJcEH1ZaIZhcFNRG9X27SSpoMNQLtSasxFEzin/Kas
Y3VVV7WrjDB1iAy6Lw93ZEBC77LWDbjeTkRFF9I8uGC4eka2wPm8C6+w/zf0zRdWoKfeRpnt3WH7
5KhXoTZ6SP79YddSAMobjBYt696OBnfeT7oV5GATur9s+NQTLrHdOFTed8S6rOwEIWIf+Jaf+d0g
JNREeBTjcDBVcNbW/Nawo8M4JYM6oeF35tYgwhzPjx339HnxjJPCUbr53BhKkkh9uPD+qJoj+/+e
kvcWNa3Ih2GGZMVahab34bp/nXDJuzg7lR0ry2O3mGyBko79d0jtifZQmLCoJjns9Hrr7bOVDUVf
lWTyp4NSOzDlfS359Jwf9qCITgPkwGvT6yZLBn7suptIsWINOsu0rI1AsXPhwQsjwdEvfr2HwhTV
fPPVBW0B5x6ne7BsxlAyb1l9650kuKA77cJYWZgNYw1k8ELF5TRU/cmNIz2OheWLBE4JsY3z98SL
h4Y/Sl+q5DmTomkp4vAJ7JMs/DUrhql3QATLiClZwJBvekFMStmkWkDz+ww8RjEnA0GE6oP5qo+8
hNG4sFMYthZkXtYt4W6wHXLynkBJiYp/BTKBg/RetqGvyhgrU65PKYXZMpbm0tiwrVtvjzAQMpxX
qyQ6VwDgcLWtUbu125WpaayjapaPsn7/4QtmSxdd7ONwb7l9tfd0OssVN6RjHgJra4swuYETlxmA
rULXtEROfswI55xc8hW8j2BtA9kK64hPhBszETEA2FT4YgZf83oFYch71FS5mSlnot/m4Jn5ShGS
MBw5oe+8b6/5cKMSfVKiH8pMB+dd7JDJP3bT2RTpNmG3jynoxXsSZyb0T/LQxKJpJRhN9fTLKHjj
VdGFVTwdk6T7BCkkry0g1fJ24zIR32yGY9EPZqJuCo28x1cdhU9NKRZkelgTZIffOsnsZ2I90aaV
DADa5IkV2P0gyjUIHzqNbXJs8S5UJaaN3ZmxtKbfhOOdtkdN4+cUVMzz/K7gb6xw+ziLpyoEVlnb
jHSsi+29bZYHMluezjar6DhO/+LEbkPRd4DnZ1omqo4suatRrtc34TCvKA5vuSauWLj2tvIC0qxx
WEyESFLnKwEhEZCGt7uSAhjeCCN+bBmQsHSWBUDYNSJarO4ts4PnhNJS3lbPsapMal7YRC7BSY5l
oaLCysw6rpwCBGhicjqK8fZA7uZydLhFL/kQModA6WRBq7Ce9kXxWRTsQTFZzQg1bGrAnSyfumha
4ZZhxLK3JcZcRsyLD+9oqp84/uV7govFp3Ghbv8NgMuNICz5/L64J3YKShtVnf9JqN4Wsxi775MI
DPH4slDS09s5+xGEK2g36JNubjE7FpbYVMxtWOEqdYCAGRSDSsFJR4TScPQ4q7KXMdq8Iz+OyexN
Fa1Woci9NbtiK2xGUq3jJtS3mFs28GyeC2vw0iAUWXxVqzh5IqtI0LWj2Um03SrOmF/Mv7brunxP
FzTKlnN7NzrTC9ZXs82dwuaaBwaXd+T5BriQFL9xBt1p0NaLV+WFbVGZjAUoIkg8ZP9gZG1foHgS
jscZSPgghzgetMQXExr+jJYzoUUYpl/kS4CZB/4ztqkV2rtXh31eatcjppDXrQwINBni7WzJIkpT
5vsMX07uY19C289ezwinhhSAcgVo7Skqr2soLnNVQgkqPSnMHa/ythDSVZm80Mgasa+7ofrJ2qJB
q0FmKJxpHity8hSox3CpqzCSLhNDYM+gg1dqH98+4R29YAaT693aQFHMBF0tcFSMvkqIhSyS2EEh
kMieynKosCLIIY22rEwNRhGp/Zmg8DS5lvJBhAn9+g1efX8820mE1YxUNbcKKdQ7pta/iXcscP0O
h1ZwGnCmP9hebae2T2J0dmMqU3G5jPd+RQ2Zy9rW3xsZ38IdifN03fwcU2WWJ/FuZpJalnifb5sd
twywmvnuwBsFjtzM881U1IqtSaxQSjp2lU+kc9yIzqvBvUg91hZi0TDTYTtBtWKBI+ujvubOBfOX
JJFKNn+uK1EN+l9YCva7e74SVyYkC7IvverXK6GaGJiF9ycgieesNM97aXksFq76Y3hM2WtZMqhi
HBpHT8g4Ic7zrNmFBjowDSOIHhTKFmn0g06eodj58asaNElcRsiFws54mvzxqFnAtkCqI1P24Jsy
iGCyl0Bd7FE3tK//jAdpsnlxdZlzKlleDNpr5tdn1FQH/SInq/8+uHznQfYeoBSPQTH+D/uehuHz
LLu9rulWjUj9w9kWdsSYb28UYX8TwrNRTSe0aBSVEvmQ8cqz4e4V82FFgEuWsQ548eIjOquO2Ai7
jquZrascu0xz8AWFc8t774idqkehN56LfCPpCYKGCWlmOEo96vSiCjK5JFZxxEO6f6xmBpCLPrAL
SO2GW9JGlA5ozYXZT8XcaYs5Dq8D1YM5aLiq21cF7sP5NJHD8ar1aN/k1E/U5HKt6/LEgH8NrpPN
c1l5rhjhlmXoLoU25/CTv5yb6RLjUiQSilbklavNwV2+TuqEH7uQMj+rJ03Y02R1nt2A399l8DDA
nsQVpLfJ6Ggl5JPEevOHsowste7cFvRE1dn4GmF2mbEBk9nN0VoeCqDgdU32XMDqxH0r3iSlFxQS
+UDzGx5uk1sw+pAVcjGekYBbNRAeukZ+GSKgyaszrC7JMGG5O0fcn6mHB78rgYY4cs51X1qaIbyB
qMnPmEwmF0gxYz1jgB+wQ9IOrm7KcM91hehhl95aBWtXZtDACglhHW5ugW+iiXC2Gfi8+1drE+hs
PmJ7vF2eoz8iVPVrh6bDVLj+wa1WL35+6o0McWWSvvW6APvpopIEEjEhjPG8AYLE2aeEun7+/04B
k7hgtHlEaGowsiq7aVPAJPR9Bx7iAF39/Z0aSEp+dLLoJkf/bdhBjlRqyYB0nKgaVmxU6y+xhcMx
Qmi/eTStYCr/l/d9GaB5f0MZXaesbUJbqtJP0hQzQOHBbmxI53icOc0wguTJGy/tQ41wZGnNTLAP
F8tmKTK1eBhwO0rW7/DfYqDuHQZU46USQYiH1TUQIRApPq3TtGwJkDuZpHbg3xGB+J6hkp1LVK/P
m9a/zABntvJ+hZ0XBBh8O+nW7/ZR0KHG4260Fod94SYXnGb/rFOTfkW2HxYct1itnHm2Wz7znxP4
S007sN2YrFO+FQ2iah7Gsu0I1pW3yBWbgrdWT9yxJz5kTXFHu9KGjK/uCH/v1zv579GkfEecJKYj
gEIXoUX/wakPQyVRKvuy0xpLMkUvoLv4W+Rl0YZapKGuwMUMq031Y++ZTxNQxcVZTqwgYGM+dxLC
XNKLqeWuakVNQJpDAhLs76GYWhOgvitnqTrxvJ+zQWqXeFHKstmGxPxA1TltBaLloRPk8/jmLgme
+xMLAenoGJIPt7BbGYXvrv5S5zE9aNGnvwjtlTIQLo4fJU9t56woFdaI1mbhjFqmgkzVMZoA8SvS
Ls34WbH/L7n9mTNTdXYWBy8IAHjfBEysBmRzy8OjcHll1A5g6iRfUpaVtOAcyLnLUaWh5KNuJXoa
poFvzoQIO06ZGVsmvuP7+Gnr6AIq9Pjj4UV3D+j8n39ywz+zOXJ4mQK/dpwKqGd6v6axbUDo301q
Wa3L2EohRiGWMZKlvVy0cY+t2xoUteIMJCfk6oCrTlzKPHLZcHJm6j7DlquW6KsA9+Rqr9Xmm0xT
L/S29OP8Sr5Jt+8umLvzccZAkCOuB6M589C4ts1T3ypwVVg5GgTy+5PPtZeqJcrmEo1rn6l4zUJB
xP6rkJVCaWuhqsj3MM/ZIBDTGUNJs0pWHTma/pd5Kk7I2agKgaZEAsMIjAvhxCaMToCm1ARHlk9I
NZHrA885bWmmSvjG8y/WV1YNNtpJZYcMAbh6vYG+3AifLBSbyPILYOBpcX9Y4TAZnVfmcUr7tY37
RWbfXa/OqLBdUO8RHk4uELdpx0PU2N619O8yzCgx/Ltw1NzPSK2L73uU2IQ7zZEDpaG0iBFppjTU
72eZTg++Abl4NxkcLNneD8BsbtnF2WXxL0ho1pDp2vINEJCtcjFI2UAt1gW78WkSxQq6lVUChBT5
dcIQVfgHNJZFToiIU6o0m0kNIDt90RH+4D+7ztvsLe7IlkCaP5kWwHSloQbEzvsA4CWaAd4oCRwG
C6cNTdg8oL2q/ushxcPS1GLS1lhw2KDgj+aZQjhmz0VpksMJ9217fkuJ0DV9zDY2XAYjlMIVHgFa
q/T4J4ke6+mXJ9/y1IqwYMkRui4eR/RJbmQbufqBxLnetDYmja+U76SUxthHj/+kTTSIZffL55l4
yO79QscNYItBz0MaWKOaf+fm0x12rKhI4opds5cCmCIXrXj4N4gMqrtrblKpKmBzxM/qun2845M9
/huMKGfNBZ8fBpCNW+arGPvZo2wZOnoevYa4b6o5j6HIWWQZRs280wy3Krh5Y8FDLqLlkECt6PUz
xwVuxaRNE5j/kyAmJIaorcT8FoiCGjmrvztHykuREJmrmd20xr7+8M5PKKjYJHQ5PQDTQkzXvRfb
XraMkbNIl61D0TsxkanRZ2Zj8D7JbsDrkrtTGoYu3q1+Fa8hoJpwYpEZb/c+HuRQu9nsjhrW1bG7
AGystuSTt+1ibldO3EDGZIbw4nUd64h48MkmLvlJX0bwHXFKdV7u5k3iw3KtLHvxAhMpvVVlbE1s
aBbIWcSS2CuXJcghBz9B5o9xVe+tUWz1dAWV2qAhBMh4pvdKHZf0Pd0FedfP8SNqKbfr8OOryKct
6M/02AwjCiS8xKYxQ1I9UAmLsu5OULiKsV9eK1wSaG8yHbJoMlweX9+Rr0v4N4p7pgjKa/SNVmq2
La2cLwKByAJMgU6AtUs6KrTmBSKIadZfQUzyYJ+UPjeVpjlrW84ypBTuy8Gd+VlZ5b9EtnQhWc9S
CCiGjaVKTQSLGiILHxnCO7ICck/IFy1AMJB2TR1ZilMi3E/ki5hSvn6gNoUC6CnGYPPec2gSOKrj
e0sKlpkjK5Gpx0wO2RJl4O6zZLFPs2wrRf9EwVn+dWJX8OHbHVAzty2af+qYyk+oQ2nYy2iCATNz
Hc2LKtxeb8pjJQ0KHgL/Qf0bQUK7DlRJwNYxdZTuAvS8tRwIqYJ1lV6U5xpYjW9cngy61TvAh+Gt
xCYFBJzVkJtYtRWT5LM599XSau7uYY8OSWA75hZ0FqtT6btNr85SicY4nQa5JTvOwbhuvn7+f4dq
ZE+9iTFEUv8M/gt2TnBKKaXfLrQX9bfC1n2XDUnNmvRk3ya7RAVlUH9B4q5SjXD3BNvgCVBK3jUL
CEISmJgK1MbHGqEhJQ/kt7ozWQxoNCSn/oaSOaQQbzv9J1iL8soXx9m/9pD+f0iLBPxVtBKxASi/
lMddCixkUb9DT/P3VKgzd3G0GsWjycT7FO7PAoe+riGzheMAyrZhJm/CZDGAVlnJEQHUyHN6Qrdo
XR9FzOROIownl8cmx8gB0FCBt3QqLv2ZMxfRBDSN7KJfis8AigK/mtrAbSj6tqExHx842Pmyt5GY
wI9M1TZqXYofqnywR3FhzHjCR/x0yYk5V0s21mrVqJmGUQU18KrsDNLVrp0oeymF1hb1VaZpFvip
XnlDdP7KHKuwr/N8/TNFZdetDblR5aCK63Pv90ItQ0Z4gNxLbIb5oEwMSz4VaOQXplqUQrGHTGt2
7ftL7nLgh7xFUr1nSk2d8JU3+nD/Np+IyMSVxs73NqSlYI+vkuPY64rFU3tHNAQjm6kFbXvM7D8X
wlzqQ/0uhB/aIB7IwHDHZfGtw589Cj8iSctgXQK4wCd0Qln/iNcaK5P3NQxBgJXGZVKKqOgigvHY
M1UX/3fbqUPadgZYHFYKQfvyDl2+aRjcbBAIxY8dMsqmhW0H15j5b7zWC4Bs4LdAJ4s+XUc5exfK
ZnGBncv3rDlfmM1iwvOUjqmtG+9rOyUsOl6fQmErGrZ3cFTyzJIWzzRnV+ugly6wcYZdLWEzfuz7
1oLniuQ23ypGYiwHLsr8aH2RM5F7CiaZlfr225BBOtPm//G+F79/Gqf4IqihbYry6RNA3XH5QGM7
k1BOcyhu2gHXa4uRx1HPo43iwac4fGWgJ3JElrMMvFN6N63Xadph7WftR0v0Bg1fUcqRIxeFtOX2
LJdz7ScEA3pMU48/7bDGPq68kRKhb9pojyxv+M+YarE8zP0MEP1dQAF9rKMLZrwxo62uUGN8lCkM
o39E/elwJj9WvhJIwkmBs6sdksEqAoY0T8A+dFJi0cKq+34eyu8smU0IMu0BNITchyMRprK16+cw
eabMdQk+GcWfJNj4Rxn2rx/YErLYWflIh/mbSbg3MiF7je3X1VlD5Kpl0XkhpeFcGqTF++ZAGWyI
BtfhFKHx6+D9wp7qlmlIyMdG7qet8RQifmqTfd45uBtEMVswg883Tzksr2YNgSwLIlbE38zotmjs
PjsMLMScRe2qFiXxeDB0xsYND2kn1wC9iMTp9COTwAP74Z8LX6XNt1w3lkucLzxTDPebTeGShcY6
Dl2ato/oAWlJpPNHgDTP3FfKzWSNqPFbKJ+fBNOP8c4uYwYk4oxvimEtoFX0CFVfo9oS/Cwbucs5
sCOXWs3HHJamRgnkp6wItyq4KwTI5lG3ZlTGpW++t5A3MAIZH1SRyqUTX/qWBWAZJLH36aByVNRX
aFZtTyb0zKiA5+jZ74itfw9MWL4NjKtdfrUwaXteJaBorvN/MGDCVMHVwZX7ZzQ0C5JZjbgT8Ixo
e9szkYplDbMsLvati+5qskGacNEn7QCNGBlDf99TXKlWiThLKJy4cKoNqu1+SkUfDZ7xCEDOkc8m
5qWXO7bKMeg/Yyyyk47qVE9CFLkVcO0z2R0MucS14wXPSYt0/8I49XtOmSP/nkIhXhyQezyCw2L3
yqGeD8IuNRcGdexXeeYT/SXC3/NX23ZlcRAdkYQeNMQ3Gnohxg9TwQnZzjYZFoN6Z+hNlb0E1fdR
K3JTs8oFkxjHWy1LbI2lNi0Q8EtGiF2yMx5u8uwIZwnkcxAVb8Pp0gIzzUQG3sxViP5mKoXo6Hj0
eV5H/DcHup663cwsilqEWKw7nlyuanUpUcRaiYZ57junCziWMpA1FL0Vi9DuJFf3TCVvlk3yUCkO
/ijm1SfTKEwN68jzDq8IYUoMtTkqZrcHJwOdHQSfvgTRxuuZ00b8QRNr02I1UwkBz2iom3zftBbZ
+040GZ9y1Hq73BbcPs6Wixoik2LzyotyKb1mwge7nIQA9BQPlRmtStZ94xUeQ6Ux15Vyzi9Pw1nV
W1HejGRKOIc0uUUzJ01YkefNTbha9TdCNl1/nqULRu2zrhJNGv5yQjfNZFNrGCu6CNEPLmym/jQw
Bp8ED/5ifz4FswkemLM5FLf4AWUqC0ek3QMgvXJ6Dc0kAtGsQxFOUi2lCZ8y9lSznXPQvn2Zkz/k
EPLRdjk7Fn/LZ8hZG6fSQmqhbe2M4EpRK6Q09xYkWrHe8Erpea1cuaikktfuyYGnLcoEDcqO4s8Y
KcejPRMLmEM+APadjLV3yG2cQ33cSFT+MjgYIVXXDR4r0dlUPFDr/QdqAi6V3rIQRPTHPvSuqLPx
YP3vHdJrq5ApuO4lhs8cDxnDBDFqlLogbQ+FB48GTI1Gc2q9tTEaxEwqQp1DMC50PUHYL2xeuTbO
uQqDqXutd+9HBg65LJsuVNn0YUzt9hRKsxVFWGvdT2htiOmDhFc5GhKxZFf4hEEsew+lGj4MiCkI
epODH8SVW2QIXExZbFMkuxIYCxEMO+VfM46gqD1TepgFSLtXMWug0WnpiYkyIDKrkRpMVThDm+vI
OUvIVTq7d8kU7CFvRhXXZByvKEnTiwrzl7SxlK/nIbbDbojthUrMruQFbhwGuulkYSZnc5RdzrGK
/DVgKFPqm+zKnCjrDtTKx8tQWKDRl53VNvUJLB8fK2RkAFAkyVbNBHkj5nQv+ykUQAtnhyUqt3mi
mHHfQB9XOhR3yopgwIp3CCKwVBu+7/eBs5uG03adb9dal/swhMk3Z9iczCT4nKXXnpKXXwP6QiNg
1ig7gwlEma9jcaABeeGNDlTSp3VFiNSfGTgZS11OEFA5+xueNTzy5FPKlB5QWRADMlMwahxll8gt
jk8YjfDo/aGeWovQq61Ydj5ATr1+869KiQPd5hiF1lQ2DVyUBYh0xcXOBMI72GBVP1sUhYRoJMG5
7J6ZeeQJNCo+hzII1g52GCGKtVkdeXC5IXRgEdoe5EsOBj5kiL44lEJi/QiG/KrblrNdhQf8aiCA
yEdqt3fnMvhStN2bWVqzsUbWUztHIK6/rMkqOmgtAI8l/qUmi4Bl30sHcBklo3ChTRT/fKPti5D3
we2FgDtl5UhGZ96miIWSypzOrGLm8i+u+brRIFXxmoo0Hd6JIaFzKrNC8XMeLgG5WfvptgaFbBYT
MpZuQssmwgHK0KMGgl9V/mRlSDS/82IUO6bpOqwWiQJ7767f8+MeqsumCuNw8rhd79cgHWK15IpR
3SIAS85oajj+NBKzHycxn8rWUf5nP+Ntz/adhprlvlV5OznrwYAd90/YekEa3JvUJfJcKPrIS/2A
8cYd/IwDfOzkefyP20BJ5YzE/AoOaYhg+jGMHtH9DNnkuLVZ3XVL608XAsNjRbffuRTuAknVvtK3
5pbxGyhvjZQCD9P0RkxuZcw2urW0fgD5L+E9DWujgZPC1ZEranmwiF3/M0/b/GWnvu3QhlKNTwcL
uXcFLMWAxVS3d6NVKGeZ25+RZt4qeEw5Hxrw/6dwq9Fj49jso31EIAKDgbypfZc3N3dFNkVeUL59
KpZAU5h8H59brglbP1YjA8qRokXoe4Jy9Oq+MV0GJaLlexDQuXpDbUaL3mU4QVpJmRvyCgOG4fty
MgGsB6iXOy8C9eHVgQGLhpr7AN1J83XfPRbtfynHxiiLHPPTUhVHg/21pvfK8N9LEMhjzMHdQWZM
p1ill691T49xcwjEYdchBaM0PPv43/6dJ50n0rLhg8JnSCs4+66Z0x5s2bhlc8RSYNMOQdGwAWIh
qOXoBgTf14D5q8O4hyQMBGvkn4DQGx7LQoBEwJJIEzfVgVFZull0+DIz+eawOIdLgEfAKUXn4I9s
9E+42FiFk0+Is2Bdt7DOOc1CHgLb8BPZfVaUUYy89oyL39ZcYlJJIUdz3duMmtv2+F38do0Kcvj3
vDrQLMZXAdQ/R34Nu0CWO2ghtrdwcGKDCUJfqoyuT4QuzSo3EzTWsGvOFwKCl56ka/WJanYvK+0F
WJkXlqpTdGK9qIGPstFJhU9fi6BTJgrrSj4wPHXLWDQJguoysSNquwJlPbb5CBBRz9lCUYCM6APj
f+4t3OgmGgnx0MrgVGg+8pQ6F+y5ZGkmkk0PH0hRGhTAXKGPn4OlLxclLSiYM6Vhdg65HiLCyoEA
jMxmqzgjAy3z/ulADRzRq9mf4mJz5swHqWgb5j7iOQ6C3IJ2ru+O+BLLjCuO1gaD8yNMT6XjImai
TzDc/RBl4sHi1pQgOW9p6C7kENMNIZq06H3K0ikwA983S2rm2banUCxsYDNL0lMBlPf3WIeHOgE6
byKFQ2ReOMLc6hCFX187Nu69XxJ2aFyzU93THiZ7rohaKrcFVtL503dzwmpxVjNPYqgetUsFASSl
O0G+EJ8LK+QD88qn80hs2wTupbvUxOfHtKEkzV9VyorHuB4VXZn6FNHXzqY0JOMZazupXb32TQF3
4+lOsg31+GFaM1hLn6P0V0I6jZtD5TtPlP2klSMRouUCSFGOWjntR0NfKdbSt549r6Ulrh/JB5MT
Vp4CSsXVJ9zLDWJeGiXc2P/9/Z7JlUmE9AWY8RzFlvlI0Z4Y4wqdv+Fcx10k+hjEyeZ6ZXNDcAiR
RvFE6gUh4pt5F30e1TO696bUsDf4cQJ2x2o8y3RG8SywOKs6o+KbNSO7HNa29GldpqUB65uZCHlE
Nfb5p8GlsRrj/3t0+3NkoM8/fTrw90MPAqi4RRqRpD3hbO1wNPQ7nsCZcYJO3zGAWEDXwPwbg/d2
uy6FQXj5VgPHydaQRQuoj8wZk7JQcMeLXjg4iqy480X2rN7sFtfBCiJ/CpjofslrLYd6KqPII+tY
K+z3HspTAE4so2qrvCBdoJrj3+m/4gLHKqar+pl7tgDNuHkHF8274dzw20HUxoiHbz43EcJjk9b6
rc4xGKyOsOrBg8KEqW1e+Z9bsAGAuqyFuLuaS52CVYc5bVKzeAokrPcExV4VBlXSBEUqCKSOp2+M
FrKKbOF0jbeYLYSW5sK4vZBLdz2t1lKHCvXaorEEBiEOK2Rkh1uHnfKNBEgoOUECvOeDk4fHKziS
TyJuUCQvy7LFEQfoK9P0K3bqFTlQK6oyGx4pTTvahRgZpBA6Onc/QBhOm9ID6fEScPUWhaOQqrGg
ddEqHcZefRrLBmiEuudXejaCmQfURgMhCYhJ5Oqsxmls7BF3g4Oo8RRfz8HDi7QA9rMYLVpjXRtL
Tuqrw2Y5SXpBPMzNJkhYSnRtO6tAIpdo4JPRGH+ppMQH1qv2pQ3IgUJK4zrAFhCW+4oUa3QM8zWi
EPPFaSuH6DYWyCBbIbsroy03T6mL2ji17gBwMvgDrwxLJ9ausNgY8Q+d1sfsxEH4s66pXikZ6WmB
8vguaFpjE7TmxDpDGRKtnBCg2eUPFtT8BNw63lEChyn0imHCoRzuerZ3clv7QzOKyj6/Y5Zn160Z
Zj3yj81lAirpCGUAT9+es2PP/bezKYRggzdepoXDTIm+HqcQrSJcxeG5cMkfQv5pCAMbgKbJ0c6p
KRZ0lW7JL2YnHpusuC/lW4yAf330zaeOC20w7c3tViWfFp1S+C0Gv+gax7JeLqcohDuktT589s8N
rXp3RIu+9jCjfaOsq952pDAK7V1OUMeICknMiRO5nyXJ0sD6xK3bvI1Z1Bqe3LG3TX2EINd6jqii
Kdg/ZpYzfarA12q9VSy9aw8cEA2nF9zllCHQS38AzYRF4Q/bTzy2rzVanHOt8WtRN6D/Y0Ssxgfy
ABjIDY3nNx6QnGGKH9s2ylNZvVIWbF4Qd/Y/7xvEQEhWnR2eVy/CGtJV2FcoolM/mSq/Cjz90jh7
67o5RQa66n+lyEGS+5asrES0C2sRTH72AWKenTjp9tLN2RjqCuhonZtfyhKojlQBZ3yVNtswpujb
/4jVpkGsdht1QG0IllxOKhowSA3PHj7D0yArJCKD0QpWPcld/7wMz3OHGuRFBXXr6xMJnUk0fcRR
uvAhdrg1oVG/K4XXaQTWP2T9AMr1dOGuZVlCjsAOSF617h4W92p4hDLGnurbvA1+EdSb7ElM9/6+
DNpt9XqlnDehJ//NuB7+ASY89Ry7wWFf0OWsJvULoCFlYo6b3YhoxEeijH6R1VprNZFYt7gO4/BV
1xVmi19gb7skEcZN/bH1783NLG6eV1RUHBtPypco16YHYHC/tXWmznLhbg7x8jE8Whcqt45gcaNu
iDTJ7pZ4dIdmqZC/NvOqvfGuGOZuskLILDN9BYnI0mYE1iVYCWiPTiR4+GBP3+MzWoU6JxW6USM6
DU7tekhqED9kZTeB9R0HTUkxvOQx7vExxd+UgB6ZmHVsrqoflhxk/2XDEywEhRfPRdAX08X07jDQ
C17jS/Op5mIiWjbFL3zHc9cLc9vkdo1sSEE/lb8+7tHm2DGy50tpke0e6ZF7PCcd9xTVGoJL+0us
LRGazDJIWhgTl+4BpUGmCNSPwhQV2kPXRCOYLxfNQqOUY9gM56vd0qd4vRkyufu/RaeG2dpz0u10
l79vIrVqNekN9eskMP6Ud9Fr0z4z7g1qxptPTbiwngbf0zs7S2qOWDbswCU1pMmXIZbPowp8GVL4
TguqhUbu06kTVd0zW5hnsfGqO77a6SCFTU7YI63lJpBnZMkxAV7kzuSi7somCEi2IY+bYpzn9udA
h18RJXN4vfyTY7Sdh0cplXmGHwcwwn1+73AHhcDCy54AIn8EpDnJFGpSmTy6+pe6WvyxCM6od9rj
4mou18urQdPJNk716PnUvEWqnK7LqH1WPwosMqLuMIQ+wDbx8Q05jeZCWf3WnnFaUv6Xq7PhSgcY
6ohSSHfhGNgMYhydEkNB8TN1PwO0PcnfZ8kjqeYhxwZ0oiwONVthShX262VrvyEp+hN/cngdcFCP
I2nqlkQPKjmplvfFR/sACuiKbZf72Zx0kG/WZADA4dKD1lfdWVTIBP3Vk/Uy3JCyKnYD4mRhQZtO
7UScFG5+sUPivaDgy7F1uiUNAGMlkBTE5tY29VH+UWtBy2i6veNEJGZi2+rJg+Ox8BCzNtDwCvU4
nop+em4yPiiS4D6b2whNn5kt7Sd0P4mwjj2GduWi7EukomZjrERSJ0uCR/9yU/vVKs4naRk9Y1w7
CvystDzbl9tyO6YcQ4tiA00CH+rH+4Od+mtFinqX/Mllr5/tluBCNBQFtehomOLSu5WsHAayee9e
4qXCiKxOO8R8ojUCV0XwCJ7RokjqyNgQWmrJ0HMrtHMNW63Exk82qGBZjHxk/IHs0RITlh8zl8s/
B+gheGMNy67QELhbU38lNDFpxwgyI+Sr1loT+YxaQWI0b8DXrILPZ6DMnU8vCf2u3aze0U5Zo4V5
qlcraWiJkPqwUsE6ji522Uzd9dA3/PoYTtW4NAOnaTmppRaWg2AjH59O2n7s2V4RxvGTnE+aZN8n
jALA9k6yIDdSDdwlZMvzk4YCYMUcCwPFhIJceQ+ExKiSoms3U2s3HHKhsNaWoB0V3bse9S8xMn8x
/5kad4oyol88miTrr8ZVjlav4qlkAyY4o/pumJLhtf6HjWDdt3FxvPWK74iNDUfhskwCZgYE0ihN
/xWho0PP2BV5Rbm81iejCVS/BCdpdePqvpffaKST595mjiL+03PLc8UiiI31fC96oW/qgpS4bcTf
20OY+IA3tUSGqtX50+VjJqphGoUAP0pRk4jOySE/DcMGLKoJq+S1zetVqcKmy2VTaa/IXqHZuIhm
aW+k6MM40n5Mz8gxtgi+SLPcvkHFj5sn67r5TM7E2MSdsGrhTLkwaPb8mHSWZQMhSQq6CP8V79ec
qvfLejAm4lMys5strngdmcK+RFuL/uoFy19X0VWhbKHNGLdJY6QmiazCYemoDZwuP6d4UnLW2k5f
CQlbJARhkQQD4bV8u3HxzuWH2CvsFjVgqFn7zmQMRLi2zi1YSPl2mMpVXvfX4q+GMkhznOyVlXmh
54Yr9+xAZC9hUWF9mRPHvaGSX5y7wjvSNgCsEnSmm+uGiWl7vxk4YnSfOSPZn8I0raGiKmFZlTLW
wZrC76CfZLUcoOn1gArYgLI5PR9JcCdbm0NC21LfSJc1GxMv9O4RqFRipOtpr3R+k+u3Se2mRaA6
92DoDN69nk6cC2ysM7RY5VdkA7pootdWwc8Bg7KXygm0MHunyuOpYqh4PKNIxx7hiJXrOvx1eBKJ
GCjzJ/dkQ/wzfAbVsUuIHvCeIKWYdm1xyHD7Pkg98JZY2uoewo2KYV6GsaI/O0Nhf9kTLZffgtVC
i4P4EDK3Lvm+i4xUOHG7EsE91OvJL9RseeCN84UikxOBvDcQqGhjwS3xB2icQuU/EofywZk9I+NX
IYqy+6dMkNDzlbigNYLK9nJIqqDmmGXcPQVScZ6hWFDz2OFOTAJbdqpiVfWVqzhoDdhCe2MCHZql
sed5zl7YYju6lIPcewkXbksbiCiRuG9mZX8h8+ZEgBY3IHSfzNDNNNhTPRsKDY4t0c7zv06p7HR1
oT1nO7GqjA0Pu638yXyQyxCqDkOlkQT6teyQhz0C9L7z+KM7EYJ2tq6sXYohLcGSEh+ZkZ61oVT1
Mm783XQADh4wMkkzvsWGq/jul402iUSBXwMiPil+Mqs7+gM1oyAMecVreR5WEkYZ0wAPl2sDiOHx
0vQ764Xp+TAgpn1b/w+wBlbA/awMP7W5+tk5MyV7GQAxR+I6i21L/7W8Fp66LLFv2vXvBjUfarxA
Jl4pclcc/ROzfJhza1nxBAzgrQMecov6RHRi2SM0dLUuyI2VwImbwbJM47Ak2KFrKFCQwiaI2FXM
AatwnO0sgZIjEZRNo2yyd49wDUc+U4mGGgBApUprzK2ramjc9T4emlPr9f3Ts+hmpWnGACXUEeU/
ItMbhwp7sz0SBasJ/+bIpPj6Bo4wLHsBqhCYeFR2HNc4ToMtxcFZNMmRv5CuTfs+7PQWHlJJgblZ
XmiTyPwKCgY2yAJx/wUpiJbjpLBCLUmNWjcLv/9feHscmwvISHGpOnbXsyS6p8wCoXcO5stvNLuu
+xYteZ7JJCZWHCFQSTnQ8/N5GwtD2qw8NPFS6UmooMf7BIrt38xtwmEOxQsoNDlPRY5aQY+n45sl
UvORnYafs1wKdDKW1U/hDdhuklJQSjoqGavhwGRAkc/L4I7fi29R1KT3yKf2MGlWfBFE9P4zyYnl
53MYKvdJF5c/eXAyIQyRDN24q0FE4s301EwbMDPzGNQlB+XZOYwuG9+rjIDSP25Pekegr8qL1Ynr
+m9VK4MHiWroGIiEJKV9V2lgncVsUwc/FdplRIcYInZfIG9WzFkAPYfrn9DgNSLj4UwYsN9CChCm
Dylg8sfjwinVgeP41uOnDkvs6ybwFDTm0nolT+/2QDlbRCBYuyj/j9I2aimfX1zQLuWLTN499AJa
E8yxoA+tb3KaCkob2O8h5XrK5x6HoUtWrWy8OLqxFn21N7CjjOkR4jJUxDQdQPCg8SXgtPmlKN1r
/laPKioaz8TjGrJITV3loB+Jn0avp19ss1JmeLVAzm64e1yT/fFDKt7ZvKXZhcL7qZIaLW9E+7uZ
Jz1UmPLIIL0nS+XB2XPgD5k3NsJQX8LX6tE04VVCriWVhJ060SrvjPaBiSxlwtUB4sK0N2hQPp9q
bIaJUjATOuaCVeWIJeWAdwBuHyKF/ZgZCd6phY4V+/J2xsmhkt60tt5fsV5QA5kbrdF2RK/cqc1C
+wnlikVbIdS2YsOCDjhWeVFs3RwgRwINcwgdq1evnu0Z1ygR7W6BGMx7h7vEYfuxmtT8CDho9TW9
zLLH08bb74QRmdWK4Dnzg7O3vRykM00NEWgfKCARmaWNKmBTe1gAKmdyh/3C6k7vNncxGEI8j8gO
D4ATVISKjZUx0LI4HvDKJqezQ+FbwW+11m6N6RNFi5P0Nol9lfPXE82lSE0i+CECHtF09tXagtUl
9DsEc7uW+GeFwgbZR6uyu/Q28XMHfiL2CVY8+K33AX5CqBbVbxAuimBKq01PKr/RkEOp30ycBoh7
C6wdMJxPhZOQcxW2ijkVviuSA5Zq2CAIjkdPE8AkGpZu+KWD5QJ/3rZct8a86eJlwC16cX8C2Zma
SR0sCoK0SPeOESlt3cEFxMxteG+LQ8dFW5vFI4otx4zewcxGfR6h/6Q2limkXUsGgxhGWqFOwdSG
orzz4cg/anR8KQpUf1aQZYKTfrfUiLnU9Bvtv8yNwTiB+Up0EmlmLTIcYPBHNAAQPJ8rxHYxZTFr
pVpfrhpAxfMXGNchC44PMJ2cD47FajwehvtyttObhjEk+uac0sqeyXwnWACqyNXbqAC4551XXzFP
Gz1sdBe8575WqEClOFmV8mT/3fCBiIPCKbVLnRGmRhRs5+JHe5EVg6IEPK39Ltz3UvFDZ7WkW6GP
w6HwGxZwMxjd5aHEkVsq+XMPrIOCfa6ObJYwNhj83MWRcw4hszstOc16MVaQFu6Vl3Oc21GlLsKv
VTPp6FkHE55w967MNJmvdHStzkwEI/nRMJmx1XSFoRaGwRj7d7bJdEveATOr+cTe4Exx3qzjtjA1
820oxH1LKpM0D/z5em93DXIfIBCxZGN7fBnApPEq4eZWj6qRZ5n7yXx/o6oeW29UNuoaUMa4EcvR
RIwEzfEMONiC8SDHKO2K+bve6JMl8v+nJZLMZ8jGLOkyMFAupluCAkoTk4KfO65QHXyMO8DGQRxy
jL+IM3D/dLuf9PrXDTCnlz+i6/04/8C+la+oh5WgLvDzHQIY+PuCnNiaIgrQP23HCgVVtUpuWlq8
X139tik+RjSvNmI2pnVkfZfhAgAqs3SH0t1ON+WLbRd7X8r6IsJ/HOpiEQHJ6j8NImlt6Z26l04R
6+ZdfzNqF3OhaKR6IrKdNP5GsuoETmJBGfH3Gw5h78R1Uz8XHo2U+QTkVNCzLZr1j/q/C7EKUQRu
pP2O4CEe95LaVRZUxDUKF7vHG3SJK6oIYR2/qIls9u28rHJnx+eKNWTX8P0JDcb7AZtvbcdV0IQC
6d3DVCXsGHBYaynLJinQhvQqxnp0oyhOh33J+RuN46/OPVC8EZga8naZ8gxJigyWSTjyaO6KiGMI
w+D6J0vyNtKfuKRqYLBdIQRRBZ2azJo8LBVXKWir2gTMfFdQAoLaoV/LUZ0j+MzVpCpaXKOxBgNv
S6i8ShysP0tr9E1vBbRO8XWoNR/OtIrbadIUIZN4gzBlXXh4wGEaHJ+hAmqbaDkyCR1Ya/BpmLhX
ebXBfMiMQaPUVNFg1DPMbBQ10vq0kcIkM41ZwZrrCE3ICbQ6pt/D3+2eIF9T1KfZXR95Zj8Rkf8K
Xa9gHRZ7pe4adVqHLdHnmgSyqzKPq+DHgnai+9k3ZFtQDhI9zCtq31+hmRzORynYWrVdVvbK8XQC
qBKoV0zZ8iFpFY2K9nDK4k6seB/KdujZi7ypz8DJtAuzeLZc/JVR5sFDnLwB5AqF+GjW75TprhKS
XaWy+maoSLA84NQzcMD3Bu6URrONo2HGkPhHewDtgY+gF+joMsEN7sswD1QiaeF31NcGlVH6DJUc
V406MATUz1GhOPt018UttgT28DNz5IpM6qXuYiDqYRQNoNfOWocIZbTUqKoVBd+cUdtlmUgjRezw
F8F+AJO59PLejQYnzeVcwfISzcJZ8QwLGTHMWUb70h+2JmXMTXIeXN3GM99ZaQE4v0hQ7wAc1aT+
9dWn+MHSLpVaa/FB9WZeSgo0AFRXc/5M9hggyY7sbw3Dvk6Mv4xoPo7yAFJFIfFRQy/+Yj571Ja1
y+1wxDux3TCrlrzeD8gJOK53AaV6mUCb5Ffss5vsMclbG8S2bgBgxtelyxMAoVn2eEvxV5WkA52r
PVtSccgoG2JSLXzWrWlEV1vNKvUO5CT5sYpVACV6jzhnboXELkNzBQd4IfG4ozOJZD3oBRrLlQ30
j7mfkOzGAa6JVSQuXbskWTyQKzBW0kU906C6bMRtoO2jiWQ0JqGAfNPWdcJHFf0l6Wj8b3bUvy0g
ARSMFPlRdhdbjbuhOis6PHe57DSfEVcMpZZMZso2DronqTUww4InmJJBStHDfPsdT0PIG/R/CiWH
rxg1KdQcMmexoz0cyPgmc0itWjzZLlR8UCQbultp/HeG4I583UWfOTdHLakFXsBhjzk2yIbXWl5N
TtXTc2Wye9LYPVZbSrPupMhkcFaqs/QzLUkY9hU7/A2soh53Mn6lMpNdv+5SLe1jxDpD8+Dz8EQ8
4dlsxHkfVjnUkNYZplGhMmjr5hMAPa4K34PUVMvMeGPFIcT1crjhDq59/CIoebgvY7NiF6CsDxwL
mlCuxdsZtezAa00RBdYgw3UfiFdPTXmAnLhQuMsIJ9Ui1zyFAgJI3CdCQbusLc1Cx/sB09PR/5CC
8aezV5MwMMo/EiIGCWiftnsuH4rLF4943mgUVLzqW1bF3yaDcXSRrTptjPliKemDrIW+eNGQcWPN
+sicRLrJ9gQvznoNIlt2OBcTfdvFb1YPlyQkIMZ4VgUCs2jez4LtL3iX2MQXVMaGKIZ/Hgo6rgHP
xe2+6dHx84A4DDlUUbMSrWS+neAUY1QTthUxazZDsAtTDhNwTUBRckvYokT/6bWntqJNwILpZ48Q
hVYKlGHFzFwjKdAWncR46SXVpTTYk2yVrTLaBgVn6TQeSSuzYLaSgcl7aQ+XJXK5Fx+v8JpNof4R
kujRC4sr0FTEbrGmjqywwLWfI6lI15IdqWJIgAGnpJbaeQ6/JpyKKb8BvEaXFnJ8UzssuyrV54mN
W4iudTn7AbTYPz42/Ek7Z97Rgqtj/aIwLhlo2tHGIrty6TTEelH+OUx3HRmpQwotYBgTphfNr+1/
dXRGhT+Bu2LsfYBn55ZGfX7E4YE4iQAsaTB0lVVWQO2nAcsSuUv1YiDahiGR2/lY+O1wE8xULFRS
cdy9bznCVXWIPbMkeltgesFiZySWh+6OaaOef+ByRf0496j24Ogm+g1/+vt5+wJI3+YII8AIELVv
7G+4SLXDCUcTyObPfdRR5JrFpv5LIkTdCXe0degJnIIXuaudu4L2vl7GL9cjNzo5mzAr3hJo4fZx
9QLQkDOV9ax337Nt7kb0KTUIY6lxCUXpVDuTn5fJSNVkbO+QWo+xvU0gmOGopl0YlVrq48XObWCI
LNSKki3Wk7RzS/v8eYPjFCBp4/U8vsy/xmsFQuN0Z2LJZxjMCafYONbBz2Q/ceIrn/uv/XmcZbZ+
+EOHXkMQ/FzXC4F1R5CnbQI9DdVzl/DVsMhfN5k9YYmMatOyX71G/D+mfuz6bMLIwY2y0yyTAr7Y
CQ1QoEbdtbyZxoNkMvSJwPudfVA253Q15imliqoLSMJZR+MOuYNU0RpPl4G2A7WMWiwjG6fupTHn
wBSs4W9WhsfRXp8yRDd9mj0tq/cSTSySIfV35+JT7I4gDyj5NLMZjBy+ZwRfD1t7Z8/E4JdjypPm
cdUnDgeb1MrDq+yKEBwDSgqlNAvy1vX5ZjFslfA0uxvmr5o6x6sadyJJfk4fw/vHLXH196SJFwQE
WVOyfsixspYlvKSyDqSQSdlKUafWt74bxJkmM8VtpduJfWqjDVW0Z6v9WPs00gOdNqJUeYtFB/CP
AZq+9dH/x7z0Zo41Jfe6I+cYvtbBlHWZCuuyKJ9JIRpDnpcgpjueFhUNKqaIP6+OKPINsEUjoLwm
KKYARZ2bEPgLs7dAU36gTtVxI3Q6318UxL3IZleNBe4WdNWcVFy09HOMPNYS9Hi7p+Tr9qNc2Lc9
Pqvt9oxowQUFBVVAK7csiOeUR4QBUTS9exJgciAoHwBYqrrqdTHpelgf1y1JO2DbawGeKLsQRLU4
2rP/LFnzygBfEti42K8P6cRSJo2snXqA9iZDyLSxh8Yf4fiXUjMcScQcRps5ree58b3QjBoStm4R
JqcdZAp1ZRqqYCdQYdr6q6ejZ1akTyNA3X4cJ9xQJ6xobWYpxx8FLJYhZU7mRJJogpDPL0UDwpvf
p7Fse25BPvYnf3vtiUqOoJ60vFnLjPsTl041/cz42mmK1O0HLJFHBDQvWOg9ZfPaJdjGJMX2FwSs
/FxoGQd3BiWoFlw245Bf/6Z52p9EdrCIzXGXdJPycNMHnk4LmKl5K08G1gPBxW/jA0Ka2uJWsoCB
b43+yJ0g3W1rIzxbh92ye7B2t2mgbSrt0oeGKlDafuM97jbN9cH8rYFMTF2PytKXnmfMpBr9aE9k
pjPfuOWIwv048X1m/c589dUK92bKaEowmtxX7r+FOhjIYVCiA8k4ea2SFkEuynk5FqnpObWq5ePe
qkXwhQDUyR7u5vlDftL5D+gkFP4lnfE0YI6oO7Cn/5Y1C2UqekZ0iq5I6SuAtUQtJnUNXE+pStTo
w986TVhhzUf2InVh/IDoJJGcM/3KirgcmM0oADy0HQPacWf7uPKNLRCao2BfNPUaOMBlNReQA8pE
j1Y+bI8WzzlY8REX5rkM+yGibqRaFMY/V+d0F/+3PDQZ/IYATGUdRsrYFkXsHkamuhOskX97io2a
6ZiT+kG9eYtH8Ehtrfqk+WmF2ZSJ9pZ42h/j3GfQaqTfAgOT/pyrcPmcmSDSIAJlrx24sYnr82k9
8ja+PMvcUE++L2+7SIZmV39bTr6hSUCpkKRXh0/msoXrEXqFmtCkB1AkJJbCQ4142LoVv3E1umYd
lvUbPv6cb3ZomwJXd2A+CUgT2jTisXEsx3++e53/a3jlSdqUbXQmZ//oaNmDsJ8zqyJikl/ORKSt
lZfQv3x6zuMyHhYgIcSKCc2D+0G5tclRJYL7YSvkcTFGh8V7o6XlJja3wBl1rxAlkUR9Aa4bZ+Sc
dgUcSH+8PGNXtHgGqSi73QoVmecTmD0VnQrhEzNBB1JsBz7tXj6VP4gCt3xOc5z2ZFUK5R6qnisL
RrK8mvtXMcii8v5L3gONVFgaibFUOBzn1+WtHxJGnenR7KucO9AsqOrul+A+Nu/2e26hrtlxma9t
jTTKhq6g5LoRQuplrpdO2RkHboUCFcl6f7Ats74O0iqTX+DLOdNiye/2tD741E63lzlyeoMTrtuw
Ug9550n/MLwyWUhm5TGCZWaatuQkKx0x3FGr25uuy7QTrqqsGOSGCcIKgxr7DAknj7yvW86QsqoY
Za4lCQEqPQt+L06jUNljvSEf52uq7Bgx6JHtchYo7EiByr2vRP4VP/pnN3EPigmwGwGVL8ANKChL
3LV7SOAQUQnCk2BmjtOMNTAtlbC9IpHtghr3BH3lVgkDEMPxfRa/u3Z35kdJIAxvPqC9CdSzOkms
3Sd6E68tMaNS/6X7eamZl+wsPUmz/1w78Cg85KlqTvRCR6vFNiCn5MaTWEHsS34FOSSOCrJAm5da
858/dqk0oaCVN8yREOWaTdwiGLlfID0Ot7TDVWepiA88ld3ce4hOFiyqODM73xKK7CB9pg7I1lXL
GY/rlkMKgguZeGAK1o1vePPlaMTSDJwNPSIHwKEwEBX52UE4ZYbqg31yBaYRde1HzDNinCSGoUPt
nk5A0RRr8lZY7axBRgEZzDRlc/I+yveTjqncItO8KwWjxTn0KgeS/1JDZ7PyzcXZUb9b9swUk37E
kyEmN8/G+MQ8hIQimxYw89igpQwAksGp3Dc+Z6nHoDNPh2nb7b5TBnFOUSMVlqPKTIUFBmW0utyT
uehzbKv6gla8F54Es8iDxQZ3Arj4rFolD1lxj4Lwg3b4enBlVlMaFykRx7OT7Vsf8q6a2qlpzvHr
cWuPFGKRdUj8zGwNVDlXHzLGES8mLkXN0fEPrwX2I3FPgQHl5WXKxdX30kNdHLU13sgGkETf5fZ+
jugSQH/rjf4dTRH2U8fPTNjRiFTF0vMW0Y2WQumKj0Vh6d/GMynSmPk41tIvkDWCY8nOZwcC4iob
KWtipeTcfxrPsCSItYRq/ZvYq2PKaAj8lHqitVQRPddVH0cu9dBGOa+TmtfJMiiH1a5vKxL28rqM
JTN7r/3LY1312RmwoeSsIxPLsMNWwg45q8t7lTzFSKlwrpyWJ/fmiBele01Qwq347oFK4rXrHvNQ
FYKBn/YBmlGcYjd7SlhWocg0PRBepRXMAJkgT6RocPG9VEI/gkOBksIvTDZDfMZlgBnn7xfvGPMl
mTlg49VXwasNWohEb1ixDGwMl0aPtiOAW6rlfw4i5KZnQ6yLJtswcJFKBZraqJLADSKtorTAMr97
I/ixhevcfQ2PXQeyOdLz/AVMMXJIhmosqhpy6ncQZjuzhtCLMeFnZJRQShUyIMfojdDdOm8DdeYr
Vjc95sHldQjb9+hRzpP29sIF1hTAPdpkvAcokUfnEeVkp5ZjvQYKmrvWPyhgj6n4Dpy7jzpLIbMa
P2XGvbMus4APZrkmR/PM+RmaCAM8SmBBKET1tIzxJBxKl61UqOMxo1/jBhJaBtBjPmpL2VBE7eFE
dkqyfiAqkQw6Ly7rjDpB8uUt/P6AXnko9TBtY4qxmQa6PdOXWJsnLbTc12q5mEraO9bQrT11J6Rt
p6rlWRf/VRwi87MCRagPWK+p3ulP03q2HuvGIgZQi3Fb6CGcDtyQPEeDwjQeIwl5QTZZGk+2TYw5
/ugiWJjHXzDiN/8lzzoXRwL5BRaZHViqtdqXenY0/rrRBEI9uwA0bpBDv6uWSUnnrsoaEyfoHH7d
scPx2HzhZmlcAHSY9CPMh4JlcHAmapA/Qn+RvVAdPdksmt+NQwKbK4rfv8M54IbTpU/U1dLX6sJq
nI/6mqbXuyZdroUjcPmNv2EMaSuQM/qI5JbVmjVliexSdojRIzUB8ssNb/2dx2UuCeNtJrT46u9s
ZFA4+HGqQWgUMERoa6itDw7ibRm5Gv6hUEXnmMkfrsyYy47+AO2W0ZTD82xPsGF9RLTA/1k+6K6s
nC3OrSzTP3xVFyMKwZgfgfDTeBn9d6HnIrhXJYek8xrrOJYln4dyY7/XkYCwMDkB3zUCpcag7KdM
HHUmpwt7PnNcGxTolc0yocFWK9bnTwYvKSvwUVGDWnflAXkMjAyr64kvxG/83HNpPNQW5YWHAzxy
GnNug4zZ5v828WHUGxdIEhEX3AH4v3UzzILZ6cAJ3jPC57xK4tp1NoU1VW1WWJBu214/27BRUSEg
L06y22eTEEAHVZNsuiggDXmK2BrsuSZ7XTCKE06jxajZMRbu6aZEnVSKr/SzWkeshV2d/5Hg4GFj
o9IaB6uQNnLUVcroCHNPDFTycpiz0chU9bcHrphXg5tYFF24nq4g5jrFXl1ofdVhTRjn4Vtp5ORx
QB8qb4idxhBs8HBdTrBD+fn7J/V3rcAccpN6Oz0XwBG+Lij4pfjXJKMa8I60fD/+RQb+r17vbRoS
oc+wLiv0UVc7n0kwfAnrO5j8WnoKSpTGhRiZ40G9pn6Wu0QD3wIO7qhg4gEIXR1uDtwJs3RNR/we
3rCb4mAhdHBs/skjNiDq/SHc0pECpH3UiTkfIIXGL4hxA4snVJo+2HSbkEqylg759wUse6QxVxMe
9sUtcWvMeBwb/dA7DFarvQICB2RJX+vTLBM4vOcEaDgaPuVnWBTGy8TAGovwLZKCCMty0p4xdIqP
abKFbj4YIV+n4RkTXEQma5UVcIUn0xtFCPAE0RyQLo6T9rijxYXQP6eDy+2XQcOXBN+ngqsaj92C
JqP0eKYMG88mQ42VL3n+jvqs8HdfpsDJmh2Updr84m4NN4iD7tNWfYqVEFHiaaFN/Yy9XxqycdTw
0I51TmYDYBNtMNQRChKZ63PxTriL0uMhJD8xsktq9Mk97yiAZ7LqBjQ2VrJg+uuVE+Vl2Br+7RC9
zEvsAHOHp1z9DkQTiX5J2EFg8Ul0M5XnvuczijLuIEfn5n5m9ezl8gBZBHRkpgTTjAat6scjiRU2
LaVOfJODc628FrQ7ImQemBYhSS24y8+eKD5HYN0ylDddsO+SZPEFFrsyg69rjljEL21rqk+rovNR
dAp18oA6cypxinfWy6fGebwQey4vuorgA9t0kWIHvQZsJNHt1b8OJTtLs12r5QotgIXr9AGpnOc+
ho4rjetMt82SIUlFtk/YWit7kI80Go0/4j12eMRia5OJEylAjp67i2cfMPkp7Nh2DAQ9HABP9mR+
9CLEZV2hN/bkbp9hqEqiRGq8qvhJgHeSY+rcla5kulGVp1xsDz/Ukhl9CCBNLcufFEYtIa0sKRLg
i6f2wHHDVNCR1/2y28cjRBOYTYCuWPUm3TUsA7akNKPf0pftRFi6eDSymSoNG8T64sgjANGpnxI6
5AVTenBSNVvYvLPxVDRUSUKFRyvQSPY1ChXammyxUv744J8SS5BcC2o8RRN/mdFHpVgd+iZIg5zw
o1uY65tDR+yDD91/iD1jE/B9z1sxVYmK5xHdXAbzzoNYipu/j9U3F/JZx8VQjZJIg7N7l6zzEvr7
kdQfNOgVvJwYmIMUht/X1wUYfQ3+16PyVgGA2+iNMQUqhsEVwfDp4NE1ICT8ZIbj0wSS6fl1Rh3a
UH5vYP6bIldDbG8T7VuWdL/dKkdnnSkfyIM/bO11NPqpPXtpM1ErU5vWmE71KS5plixXJQo3ibXT
aTTB6CPQ8KU+QiW5R4PkEs//Gyrigv5dR/bgK+0/2unAhxFyXF4y9b2LT7W8qfr81M2XnlAaGLTX
95ls8Cjg3cj/+1QsGRdFavzC0PhZZy2L3lVN7tPE9FKbPuVJO5IXKKw2X6bN08iU5G1/MRC9mPH7
1aUBYzkcN24YVTQEJGu7M2kxDhqf9PGQJ8ejGC0wjuFczaMg7+3l+ovMr/jpqvLkKhHLvDmb9n4w
QfUHSW7aIXtXcrSrun2s6eKNprmLA440dJFmDvJzYk/lFvzYFVC50kUCm328h/la2wEhsc/lTzF0
a6ObL+moR+9xXRI17nv1PffiTJXqptlNoyYsLfnhdKbmsq5axebEZHors6L9rC942owQ0aXJPOXe
LXBN1Cu7l7Yqk7/1aS5O8ZIjPvv4NzfFtmzdjZv81bBEjvbtTrBf2Ff7BY9D+70xjGhz0xt9Nc7L
zjrqLloL2HxqmHjeSZh9Kcuy3peKuqjZ36z7J77sklPlhS+LIHVnNLWZmWZPGdY2N+8OG1tUQ1CA
65RcP11AzkG45t3GAp3uvf1C/rEiF8Q2h76Hr4d4LBCCa22HA9XqIwQ7ExSTxsiii/KR5GiWyn71
u39ImrZ4nm2/ZAWVAlcNmewJl9GmM7mBqnRVqWQJP6eGTON2juJDpF7l7d0L2FuLVVGHxj9P+gKC
0kKKqK2HKMtXyVxSRgmA+klFPLTmsq1WwuXQcQ2JAku6lOHcyBGVYADE7y3hAy4LH26lCFV7p7aX
hFXnVop+MD+YIsUlybOlcYYQsjV0H/7oCUdWOa/z/RtKlq/ZCsyoYppxqSHIimYG8AMCN0Rc8tVK
e7X8EoTXSPfHXuhwm4CQGeqits2wmLa3tpAbAZbGHh9KFJtxqtvznjOq39nvyJ3Y+uBlGoibHBAX
aS6N70MyEL/DmBZD5bizEEwa6sYQXgCLyAaNr95wMyXSclO85ef375F1zbUggo+wmprJB2l7/ug3
ikqj+Jr1FouGXB5R4yFrXJmRHaFQuj4D4x2675BBnOcAy04MGCo5r5UU/77YwatGe4gdDfJmEYBc
t0Gcv6ucXZg56gtlC9nm6FqjfCnC6QVv9uofOp179sNAF/sqkbum6r5rF62cDy9hG8OPUfanZP41
RznK2I5wUmLw4blkD2qZiGyDSup4X7mq9ArNF0KaJ1ECim073IyzvqC5ff5k650gt0Q6fKyuhnb1
kEOS+mt4oUP77IS2+DlyHz7/ZvVxpSa9SUcZPTVBppvFKCvBQWOB1jSnF9VFj51CkCDP1LL4XKkX
0QqHLMXrEDO/VlXZVbMGFvP213Hr95Ky8kRAKzfWzGdknEireGh1oFLZ+cS6xH8YDJWxtoyeEIk+
olKYoBgBgcxSzWW2AUDAVnVT7F4XAi8ac0UktZVvwOjGbgvmDZnOsrzMNKZ/1f5vS0FbXTWPDxHg
KV6MrxDFyoQb0IaqWoUrXeoHMYDhQv6l27xyMAPjFJ/ySnNk84WSygRlh+y2ezrj0LJayRxV3zpy
furOC9qvlsMoPm38LtaM8ZnkAQS/kx1El4LadIgX5JIIlWvdKtwFl91sB6wRdoF3Z95oyPXZ6Nn2
0DeNm1lbU9BQj8Q9OhoBwAEQlnQfcxyulbuVbGv2b6H5hTu8Ee0CygDaVwj3zz3ktc/JDpnj2xYU
gt0OtdixvcGpIq4WxLSwZkbIdjlVWybDTe27UJgNKOpa7EG3r10t6HklPO+ZWa5N8Gz/Cklbf8aV
fGfG8+BSecMQtDy37t26xs+rHG2p3KB9nR+EjYQ48fk5jIYi+GerGf9PM2m1wP9cjjbYS/4XVA6T
psboaQmX0zG+nRWnua8IMjvt5nVqh4zatHpOt/9VApRlb8dOLHHw7rQRefS+QKB/Uazf4pZnOdSw
4vGH0UqYtbdap4C7qJRDsY/S7zAt33xisWw3XUuP65Zk6RbduoZHfGoIFRzY9YeKwinLggjiH31Y
cIzreL78bsneZBsoXbvwFPwg9KiUeX6C+bB3n7DL2+yPU9r46/XsAqYHxs7aojAUKHO3qjvMk5l3
g85BzotJS8lU3P10u+ScoL7cjafwrzzXQnxf9aNvPApM5RCmOKkCvvVZ7CLJMpGaijmF9PPSojrx
N9ji0gT4ZifefH4tkOYTbH3Rui+C51+aFunzsdjRhXPIlVgM95lWZIAgKhfsRAyZXkYmo6exyKlj
iH5uxv/vvFNe8mpxEXyAgv13iVS2zV1IRvPSxHFCgx9KH2yPvp3A01HJIqdac3bMbDgkzwWBJTBz
wQmI+9hMqcptHjpJjK/0ZcKDkmFCaAp1WnnwExBHXwHw0s2H/MSmdQaNc7NWT62l8Ja2paEu53VI
bNzzM1kPG+z+elb/50UcLBe5k8m3RipNxsvo+Oc8d3Zq9BSVQHESoFJVBvGnrsa+t2tCfqSQkM6X
rqx8OvshOm58NQOOICyazjY1B+eHgcGlxD0QRm9zkYtNIQW1fIt+Ahr/6V6eGWJwUboZkU3raD6Q
SJ4tQGr4ejm432F/IRnRFgdDnJ3JTOeNXs+3fALAIHXSUQCYX5f+vfNM/vN8vl91u5gUTIg4snX1
Q5RqfwGGarGjTdksZbv2Uqwv9X1FON1l7iET43I92lEJk1dpHXBDDzwvMr0t1S56htu71W5Glh6G
W0EFQGpyTIcmPkddCS1/uyLcegMXh2fr0fxSbqjlJwophw33c4zy5cJ9ynjGSsM94m/UAshJEjFM
V2MDOwLnFp6OzH8UcAS/hp+REZNgUaOCb/ocfhOgERNyJ3H2kylDt8D4msgptQJYhkFNdjcD7nvd
200d0aDzL2FHU0NwYwfvDn6i2As4vrzRz8LHCK2APZmf7QLYRpxdUTlFVPB+KVfLjB+jCWAYLRsX
wYAhrIat4OZJSvUU1DGrwSqqrpAPGcXg8EuOxp/ZJ1aZ9r0OyEnOukKBjDOV2Pf1xSfXNkLkm+94
VT3kiab6/Ax8HISdY1kZAOczH2VgDvLyWK/ggcXLLmpqD1WXdanqGPt/f6qu7FdcnWge/IH17tPw
WvwjG+eQKlL0AXEwL3jZVhWnBYVUh4Q9xVPXNu1hQ/CHTcEkhdibj89Ejq0mmNHIWnG2Zx2tMU/L
IRh9RATyUIYUYFyynrvLrQuKoftknPVMeV/0gu7Qs4xmd+2GfD9phsEbAI8uEYjYzC1IYsjQUON4
x0IUHojbkihvslF1hlkfCvgxJBOli/qral01yNpqL4GzmL3lHh2Dgnvs0wDHsWD693kIIkri+uhC
GR3mRPR4f0/cYKgi8JKyJDQyuJpyVj7n0WplvFkzRde4QHokBXt4Ak/coaPYqYxS+1pZm2mhocG2
Ii0BlAgwMxivCWWhQiD3JhnqL3ddfCwZni0aP+HLiIGI1YERktsSGDqhQLNQhJ7q5Gu5+JljOWT3
vFLhM9S4GJ0zaCes7Krr1CxbTMbPFO3RmxQ4zT7WM6cyQ19qvw7uME8wmlp7kWuMeZAt7LLsRG2Y
rPReKQK25E4S3o0LL611JGQi/6K+wtCnjXlUcWmR9kVQRxGDhqeSjOm3EsirmbYInz7RcPBZsuBV
7KYWILVceqHVIkm/+rALJUGqWTj8w8hCNAteUTOXMRNmg2FfqMj4zmWIUuyIGvi9f/4jcYuFFB2W
u5qBko6vYfz2I8bNngoaos1MQn0rfFILNHrQ/tW6YGhFK6TgnmmRBN+b/uvqUsFbljcwmpmfmrU0
8SVTbKrXyXXYX7DTa023k2wlDeWt/t7BEVDm6HG/mUpt8Idq6QOWDoX8eARswKxCzkfzO9eZ7SW6
7x7eD1IlgpP62TZvLWP/JrqnfahERMU4G9uQS6NpnVNteqjoiWO0RoOqEjvndAZ4vYTEVQwKX9Nr
UFbTevHcpNQhRjj2w9avIqZjtYImb004CMVdpe8M59J42FGDSnDEClcSCfhI8ZyOwYqYSSHe0ny0
QneExzjOB7+ZPi9mQtzXmt9JOPClhpCfQ7VkyELDWRCydZsm3OTy8WEufa0kQcNH9YTl3yQdDQH/
pGhbRB69Q5019q9R3z3nT2GHU24zYWfjQjX6J8dXSSVVo9BjfFNXy7vXZ5pXDZ7/voBTTGaQqLu5
N6gI7f7S4LwKiGaK6LhNlCagHtbXDrqqElYxFJnM5na8xSHGty2UzfmUqonytoMl6bgJyjENotrd
WtPtLXfnT6h49oTrv3cbLILgli0Wsldrfoxm9b1RVH8gms2ccgaMzGf24cx74xSlGzShKF0Gp023
sQ1bUK1LwwZZRnWxd99jpCRv+zQb0SMyqDSrWW6wP5ENQ3Sdb9QO4GmfX5rnZ2HPYXugXkSBuZx/
cwQUxq2B6ovuHdpQa9IXyHX6yeKNJZ6Mn6O9LJ3azsHZPPtkVsfjt+ob5a3LP/gxQgoC1xzeDTyg
icW1mLU6e74aXqGZdZP3l67d7Z4so+AjRqjPDq9bkSusdxv5a9Tle/21DnUegt8zNtCKGM65uAGh
Ea8sWPskD9sS/rNFDjGVAwQWSoad98VDsgNWqnkjzA07LZ/hrRy2BgPbc39XgH/bwEHqP/DhMvyS
9zvLxZnneSxal0L5h6vF+uH1IMIzNiEhUi92Qmy3NmcWX3K3610zBJhY8OHVykEU+Sk6zDApMkeU
/TlB9Ujc5XUF+YUf+f/xJ70vQMFwiDKSdRIOcFzRb1bgGV3NK1N4IWc1jYaqrsMBY8YWbMqjTsB9
Uw89z/9S942PxLOC9AKveF/s5yLCw9movZUIcK4NfoCLVBRrMA+swq9DNkwURmKLJzTDWbMsxuBN
WKjWv5eGdHwWg+WsY16kQrigWHq4rUi9vUK5vyTzpChgUbWtdQGv1JlM/8wHahl9JXLTbJm7CyXO
sLtPsXmxwUhsWCaHyfwE9WlaBPoB6qx7vl3YDU11PtMd7bc2mRxRZLWLjWLc1sUqGYGnOEvlsOjX
AgQy7K38JegZG4/dYhma3vBNe0/yA53pwBOVHW5fwtHqyOBooSwqEb4DGgrBDWME6PajIcokwqc3
PVRLk6a50523uF3q2WrYu2AXUO70QfGgYT2Ngsd/XTeKbmra/LNyKpnCpmhfLOV1TnEiJVHk3YrD
O0p60fL0SNuUZAqRR0Ivrlayfn7HANPTCIwjB+B3QG5e6NlX6SFKkAkKNQJEBmAltfs9FMcavdl9
rI4CcM84kuYMuN5pr1qJXGmHiaDD+VYFDzSyCW0j2KuT2gaUtbp5QazMpgyOEhxYGUhi2pPfk9p/
Z4vt4NE9qOrNejqY6t2ICRgy6Ji1FFA9NDt76yWYNzM8pmx9czHZYf5VW/3viDeSpDbsKhAlcDC3
2LXQRE39yIRl3fAARVd0gM5Jn7v9QivAu+SVKYr2kurZ4wPVhWPOHzf22/GihuJimmcd58OJdERR
HVzE/FmyKIyYthaFD0nzEMpCJYzkT0U/fEAExLfuaOUvkSpiceNCXf2mrPdgTCiJoGaHd0p2NVmV
eiUmJWD9++KwjGbUskkfcLpeIDgZXMdk6Lh4in/fdKQrGu7DaODiXOmAeMl7DMV7aEtsVYAfDWYh
pfaKxYh0aiLqNnbIvljtRa6q+okvJBZEiIJJxbN3fPsGLFXK5/k4OjzL8OuUktGNQCifpTT8bvaY
IyrKPXlWErsFhWzKPaHpdxwqCz2hxWeOxFgp7y+H95Qke0eY969b0Eu5u0pmcACUJd+h7H10oEu3
ntcGIdauGgpsLs4LaJlYHXh79V+mVPSFHa8RShFyVbwLchjt5XhTkSoODi64UWwZTAkjSr6WrRij
bEVRkLvnmEqToKBiMGXARYBxpJ9wk4lW1weQYnSJaQ2oUcUCCIhewQGiBATh8i5GsOvGjvqOecSk
zke6X0BZsFjAbWctwfFllQb/zixLGLpgaWG681UOKMxjwNGoCfAD41D7uCdheqYN01HHiukw/VHa
ynWMhRsmCv/QAirZSew3leZqcxB3lYAa/gOCpvKSzyewgcMIbIvKuyb3Ki3eS8bAbpR6CeomcKrI
+4XrLvvEXQ3UcSki6ZrZt7T6blZglvuKdBr9xK4Dm2KbdxQSKwp5XUBJplIIdxDUG6lXipte1hCi
HPM/RPx1MzxUBuL0sZ+BmF85/vRR1RkNqzhpilHT0OTWYTni3TCvU3G68DSiUrlEqqbMkBsyGAwa
R3c6T29XZaGGO9B6i9AHe7jRYBsf0gX6xXUZ80UxE3zx9CAcAQTP3Fm9j23lPLQqaIlVTOKtqIcr
a4NaqdT/+LgTx7NeXgPBFIKtXvSZfnz+QwhAszQP/Th4hUCdI+73UbPSzS8Rvc9EdRs23SmxDFGl
pPn3Hd3KH5GDldrpxBPFa3JQHTHC0OWQUfspFGdSTkk93TNE/dPD3Vmj+E5A6ssgqdFytbjiG/Um
tTjAnMCwjHBsM1s6zkugShJOpxRJUiTckhPGZxdwRo06WXOeHTbnZWIEMj3ki4gagKdnINROUQZ9
aUiagNWE4Njl8BBE4HNC9MyjVG+klDrFYAsitouNKJDFaCfnMenlZzDc0UmBYsHj/KSaNNvzHWrh
z8ieZbckCMlR1UlbMeLamGV8pEdBP7cadC1PNx41/oMXYToGT6zXBkxMK/nyND3vhZ+Wz/GzSVYt
6iVVoekTplRGlVSLyaBJymeSuQq5lqr9GG/sjuiw78p9rFNgURV9KX/om2qDRTVz+aH+XTNE6/S6
fnHY3yVu5Eouy1LrKIY4LR+rOhCkaBFrBCD0x3LxM/vzHmsVqBHFhMJUUfzxWp4vU2oJKLXSBJl1
Yg6D0+yiocIQw+0TAcHhiiqA5V0Qd5zKruyL63y3y0hJtpaDEd3CfRNcmu+eXVN5MA+MpUk49VAW
UJjbPRVbY78HgKQlkudHgbckCnW+n3+yjSbZk2H4mCWQbNIa7YuTjuMBQd8TKcrs/rxCywFFdnrV
j00f0C66RVNQB6IcqBZ33sj8aQCGavzKJhVxBxxV8kLPJaC8uKhW98z1sbmzVU24+FJ9KYqJ+/s1
fKfO7UXO+5rBwbNx+fRu1suA9TlBawFO9jwPhXsXpYbgaiDX55c/2oQrmgmZ+wsrJXYY5iVx2yzN
ePS/rPvBDxmGVBu9gZvJ1Fi5/vHC4TYoUwXFhxIr+Y1JVIx2aITAv0Qhi5U4KUUcUkhKUlpUzz/f
Q3a1yTqL3p+d2V0O/BlE9mQFoLlYPDVa25q4oo6NJthlIX2wVEv2MHLJEpoCpRz0v8tk+O+GBYfB
PoYhBWN7oVQ1pwaXYLBGr09yZFlqEEfyS/5vIJaI4AIamOoSf1DlHRHRZwJBvx57mq4KlwmpWpGg
chuwJOHNDqfuCYUFLcoDj+GadTWKo6AxbsMZ0rlydN3lx9i5c4y3tUNOm/KkN4o+CHMRI9kPykZ4
L28drp0zedsYpdkMMecgl26Ju8dZbdRzaCK7pTn2wKNwboji4XGLf3+SoH1RD5O835PwmQK7AX8f
QMHu+f+Ni8jv6uxCGcKNcXGabxfws48csGeWtFZ8tLZ5DZz9spjJOu+4gLwAC3pESf3rNWHeoheq
c7pfq73ZAcHp0agvCh+l5sDpUNj0Zt6TtM/Muaz8zWgQS4NSgUYKyfvfPSUhZA24OcDUIZQSwayU
H4jRFmvS7iw0PW2zN3zGpXTwPdKHxPnTfZxFaEzPKNQQmpYDXalACQvXxxe0cYZFVhQU6LoOe81G
vn7jQQC9yuGRK/Hf/NfR3/26+xr+aepo+VfySJ0B7mLn70E6coH8WOPG56YIKO0cV5rxTml/RoXD
zkitEouBwmoH0LMiJw7qEl68i89rwyaIRphwdl/pj7m0paJUUSBF35AFmbdSm9mjSZA3c7zLjH8u
DPTccjcxEPGOsUsE1N7JltPXLCkeQ0GyesdPLuYMQ2Qm8vdz4v7L6Y2vWWR9s6ygx8dx2b/ISQpd
UUWS6wtmm8pArQBwJ+DeT91pb5oHAXZTxQYK46J/BqSJQ7QsgFdlNuE3zBovNV2Bv1DXcOc+HVhI
QRZJaKwbHiK6qND6xxddvXisutXd2gn2wyLMnzpRx6Tmjs4/ftp5ly6l/z4zH1X4VqKR5hHVYjLJ
EXuxtU8KBYRouP0xj/9tV2Mg+BRP+OkS0yck+nErTL3WLDsC10dmKEpAVzVdS3CqvY9dZdUREvpx
9SlWFQ7aUt+rZ4PX6QSStmmW6F1QzYhwc6MSo/37IKHHvmUqK7C0eAneRwdSx6Zgku8NF2TqKQGl
Hw81mv0f9s7yBnHP0WA9NJFnlE0oZH1KZT9qTKjdKoIDSteWrAM9Z8sB83wfalqoRf4rTVerWful
9TZgR7MveJv/CVS7lQ1ZDHKkIBhZH2Hk2xtH64ItRLdQohzMZJXVTB/Bo+sNgLZ5RdUh1EfbTSv2
lbHSHFFwWlqMXR8yUO0dLEQk0eLsKwWgGxlwhmOENrS1A/N5R7CZEGtOI1Dc+18HewFsXIGQ4/g3
7CAkb50PXE+k47V/MsQmVm6RTBIfoy3CVOZ0ZDHAeop3sjvJqy/CVoE/J/vBlssO/TJs7BKmRSsd
WEasptZo5DM+AtzufD73FtIgDXGaPkEQrr1WtQ8lG6G7zGHvF7Ga7Gr6h0pwOrt0APUHCpP4CC+R
hQVwK4+ZtKnL33kKCvRagPiHQY4D/1zxMIdiNqG4bahAVH8TBCBEmm8aTsNk/Yy+fDd1V5sTSSF3
md9LORibFHi82FczpKSM+1UY6wdmr6H1iHYaMEtp4QxO7rrM3ukYpKWopkL/jL+4N7BJu0KhprFD
8c7F3L3cXZUfQ1nr4SbH5POrwnPsIx8YeDkdWZ337GNrp6tz0XgsdUr36Q0parkBUWAWWyaogbfa
jD8/hgtzXSALFN5V2oQDvf0MgPB3JUg5zU7y7pbMzX8duciAjaWNfIQtOpDK9Wq+Uqe1WD9tZFIO
iZZf+oAztZ17fUhMRebevEEpkL26lQ+Z5XLpA/0Dc1ohJm4gEjjmgK9Bqfx6TTlR+O0rTjht0NY7
d6ADFO7D3vgjf8urAx9zp6C7jVLEONM214qba84I85rZ69s0aQRdx0FUbuYmUm9O6wqdy4GW6gMD
3NkW9yqR6QKPSDuAxYcTVBbIlciexRPWlJjeI8KiuXHHjo5Vkhlw74ett9vtR+ycS9xnq7Ly3j2i
vts78jaPuBGOR0VJGmXpE6bXSLRLjmkiGJYlXAOGxixsCIt6vxEG0AR4mZCsM1XnxM/xssRpZJQ+
GIDyKhvZkeLxoppb7FyqkP8i9ybhhbkCXFgF+wxiGbwz0XhHGX+FZ5d6lC53iNmriXSum8yXCSw7
6ZPHGGsO51Xjr4t3SUFN4RWWvVAxSVFEBgThXTdV8AM19CWkaugdqD1jSiieQxUo4Jni8TwjboHp
AgFH0xk0iz4epdvXk1zMqBCf4Ad4bMcmU7nuIW2W3UeygveLL1GKAFlYzlnQhx7mN6nrUOj3a+4y
glNRMEZzF4kmbvhocjYEJ4O/ghbPtG6ksXdqttDV0e4PAa1pGoFcAEBkVCYT8R57Zxw5o4HibJhX
VE+nTtAKzj5gUzJsndAB25Me/I8HnMlh+guUr4yrnHCaFsDMvKjckyxEL7zJD5u38NsvbsMcpQtx
icQnrebyPZcq7KCHBHnPRlciSmFbPTJzpQk7sAJvWCmghhyqHkUprtV7jzSizo72gPbZCniFnPs1
5fpr2+S9G1dKeckXzLfOhrhgLto6lZszjZdccJzM2VbUleo7X7pXxLUoq5PLRFkyaOkwkTiOUmah
P23Jd8DWeyxr20iHtwgVbrZQn966+aKktQ+7xP0HQYHxK/4iyuloEZynhDCbjdkKGBUSWF+0RldY
C1ht8gU3PKQQaJDtcFiRxCLJ/N8hknusX7oNUnWV6LiHSo/mzEUxMp3Kc2heEGag0uBJO6v7nTrM
6WXBnttiz3Sg3qhxh7o7ifQPMSq02e/Gqx+ZTCC1EkrxgbQ54Qo2QDbINHxEmuUPQBjBNzKTNhZZ
l7khhlVDu56Za8ElqiYy6239VFnWJIWu3SQevG16ySdMOzobhEDv9gxM+G95J11E7meHzbJB7Z7m
EOhR1nFRHwYo30kRTXABnrqN1UVoE6P7v0bzY2coT5kMi1hiNgI1hIPqaiutzN9D3zDSl80/5SRA
xuuLGilHtDyvw171p6HK86ua8SW0LI8LzV4s/MWluK+70pJHZtcP5wAEnFph7sAfIgRSPrYvWj7+
GTjNTjx7ok1kWc4tcoGYKGAFbXTVLD3e2cXM3rYu4NcQau18Kyljcu1y0svKLAzcbqNe7VJbk2Vr
1dIULHUDvb6+FuQs9+Aue4leNZrBB6yzw1arJ2cXzV0Snxz8cDMKCxw7moChe1+1H+CxLOVlzccr
TwbmG10xkLRoBACLmFHABGLRGbdLhTVhRliS5xJrvIk7ix8tWGhhWT8yhdb+a4I/jZdpuGAeDWtk
0p5w0NMLTKYlg2CfAEqnZ2vJd2lCdQ7Lb63LIEhUXCDyPJzmMn9G0lJeyKPHlSB51PG1IsO99VMg
YIgzX1K9HP/Hrvb09lTYgNvAeY7ubn5sPomAvuQWXyDoUDkghz6qkuPZAauVwkO6k78vRslFx7Sd
M3f1KYgDYcsSWYBkcIClCqLs6yZ/t154QfM0HFAWxAlQ50cuTp2wGtQbJmD3hFveGONqn8TQb2w0
XA2Ixmgibk7/FLeKEJcpWVVDMoOboQAC4zDJq6+BYsb7C57kMAdIUXPpuwzL+qJZVaz+JDVjD0PM
F4td+nFvabxNEICL7z2E/Kp8Bc5guvDFUJTs1BdUL08WIa8ctyYE5EEk5tmiRsYY0TkdnEcjPhpz
r/uTLGrH9aP+pYgB92b8zZS2SZUfibzb3J2sRFpx0psQfry3yaU5T39p4ExXFesLiTGfMSlIlUr7
LTemCcPCMxifN0ahUeAb9sV/wSebzVbXlf1wrAXcYMT34vtXpd2/eohWaRpBg2NDHrnByq/I3SeD
5b05l7j/6QfJtPNS170J87X4LYBUuMZJej1jeOa+T/oA8JOXa9A4k51t+hrGRy3qHMs43x8aCocA
l8d+Fn5k1xmHVZl7IFU9Tcqf0Vapu/COwKYATzljhwJeUCOff+PIoqruCnZ+EgzGdpCAtXyX5L/D
NtcEGWBKKYO8tUSVBMgHcYZuy7pujnKnfQKNH+2j0xfJxPn4/OOJoAq+4JArCmVSA6twQS9egGTC
NsQcZeAyJFe8Za9ABmFsJ1ncXb8GVQj/k+qbGPL6KXKLq6CWouyCn3fyWEC6iep02SD5kQbj16fV
YGc3LrOUvNw2/9q2ynBdtHf87C9cMGfJAHlZ2X1cilGO2QqC0HZH05O7/jVyg4C3YE1c9pkqRLWu
u8JzeSwmqLe4ESsPrpLaDmCDx56MnRwPs8XtDj/UVvxfj2hyGd0DYRDa5A5pm04ayR0WK4zrwryu
AWBcwsCPC0UwB2rAZAN0XrG8mcWIyb5jn+ebWZ8LqlYsi3Xr18QZuKY2/leOK9Vu/L1P79MDd9xR
Oz/Jso3ESrRS6Bjl3rvIhZA4F+osd8Kq/OV5RkaCr+hdMu/3fcN4PjAgVG2ja+o0qke7R2W/boHQ
MpZHlm6JzfcDqO06yhhGmlzmgIwADdDFXl7gOfzz/leo2iGLvqBEIWf9NZTnlIS2t/7Vlryp4OAz
1X9bNVmiyNjz2ArjcqzrpQr/vy4NW2SbzBwigg6PlhlrU31DtSj0rFJMXEoZHMKOKtWegCWymVyd
O/IVskxzp13W5oLswRNqkzwgiogkzExZI1GdO3rD6IqLLXe6p9KUrN/wrfj5pqRiR0q8hetXxfXx
sK6fIpEaGYyotmnDc3xvasqBOXjGU/6GPFSnKXJ0LEWwgxOlcoDFx84vW2WYaOLMNciFPMX+0NFH
pA5MlNX+HKiZYR8hr00kx1yXAJngiub7uNh6gi7oYKhR14JgyqR79XuqlUlvQ9Yqp7Pxq01aWXfY
9SkuFh4ww3KC3abkxx0BKZ+ItfQ4qj+mX3OjFEQdHsvVCjCQWmneoaUsPXJ48DtYnfD/pO0kaQu7
V/EvHtXqDNXYEc6gyy/UxQngcHVqRANJ9pWhsveg5WgiOpJfQo7w2q8pxdpOTJqneYxCRpl9hGWz
4ACSzNxEivux/YcsD5SiIU0v9B3y5PPHJPlASF62rMBprp3g3BggisF/qlbPBYxYR5cT3745p1ac
Mqgd6Z5qsfucVb5E9R13Bbt80eyE+Rk1eIokC4+U6w4vlydZd1tNyIzHiz/geqvvUI1JwGmN3X5c
X+Awh+oypNMXwj0h4aNs26hKP8uwV2ajmhuF0x8raY922yRamnRu6lJp8DvSma6lvTloq5OIAUFm
SVQ/Uz7279/elPF4L4+3RX4t8Dd7FKff7yQHsTWAiJqJXciumf09v23Sjzps2oO/pzrNKb/ITlEM
qv38SMaxicNcszh+fWY2jlNcKggP56ESo98IhsuT8NvVG39jb3qYqDBX1rLlhYPEezfGnCc6rrjE
j3uCeMq5YJpXMqjiOJvm8F82tcE8irPqnOMSJQBq+FvVtQFlcvWznTfycjyC57r0OAw8Tyvcp7qr
2PPhCdiCVW9QEKHZ4R0MCOWjNN6ip0tRP+Lc/YxaTDqiWPxdAPDt0siby3i/bdPgQHhAOXFQQ5el
ldaqG38vFbYIk+HJppOoDmLuhvAZXYlWS7rutvFhc2V5UH0gWN9EUZZAnU1Oio82GI81t2Y2HFNz
YONtoktTeOiAC3wxJnVl+Pdp3Zt4fPUCCjqLdEBS3aJyUpowgSaNsbrzwYL6RDcrBdCbK0+ZPulE
rAepOYvLWVQrXhz05OkZy2hRzP/IiShxBSv/YBGuTtxVFf6BgOk3MWsNrW8FVzDxWbuw/CN4KnCF
1OYHgP0hpGwA+vvqns9FlZ+4OwgemkiFqt47hypnLzuVKtpoxIMa2AeGpg4MaU3jkcpYHxaTazLd
dyg/vmbEfwG9RfUx4+71HpIGOrLU16iVDo0k2sRmNVILNyoEb+WwwYScg8NFDlxx30fQU+MAtXh8
FHfaPNncavmlGEbxWcfNfk3J8oJlXh0GW8RMyNhEx67w1s8LM658C797B3/m7pydpxZ+xAFwB2IF
AJmyjFgZcidUtDR2JUk3fquN5tt4Cy/909EAFbqOtt6BK+3QTxfZGsDesV168aJtlDuBxui1jGcj
sRMvdveKa0XCp2TcTxTcT7wu7PiFHNZT0I/CoKL8lhsJ/qspCxG6eUQ6AQIdvRk2q3Rzm26/tFu0
FeX3NwZKOwm7k8c0YHNFYJiGH5JOX0T5sD/29naY2vEcbLSpWyVmMvq+vUQ8LpDJN63DUWohu7Mj
TaMXjfxZyerE0+p2vkyUAet5JtTH77YcxQTznibPk1gR+lacMEe3YJPHW50JrvALKwDNNCTi2QYX
d7yuFsHhMDzQKjFFTjZ4slupYpWT5SRDeUiJy2kVgouaPCxuAJu3VS/9cs9X9AIkIOhYF2SIcMBg
k5oROp0YRwvT0oJ/8HfESIipV6sHQgid0jC2Sud1ZKVef0oBK0Th/I/v2ROC+jJR+GoOlcCqGX0E
FS6xL8UEp2jevzK/WF2yt21XRSar2LFnPZ2dlDyX0LtR4QOJOHt46jJqp6zCdi6YZW+XZpriLY64
N40rBx3W9Dl+3HH/O+V8KaHqbMlYKcxLMXWjohZYiUaXj7+oYE+PjSKJm0czSLB7y8E4+ux75pIX
GicgeYJREcwM4iia1z59VkX+NkG+Gm6QmZNoTiTxhSu9BxUGmV0kjEvq1XmBSa1XhTX/v9XJZtB6
NayV5iTvBsp9d4zfU5bSUtuTWUHHo/4qKLXk7V6NC8w2XCi2D5Ytgt2hhM6wyLTP/I2mo0zwOL+R
QHK+HrvBjrTOO/14WjjgmKhdgrWURE9O4NFe1jW39mq0XwiRqVL77GklmcUPnD4CqZFhYDIdVicJ
cJwLX2HJw4csGppBwKPlLalSpnGOTEC/bOdeSF5z+tfOCAb6uBgU3kiWCpdEp0H+vMhZOA++jM3U
ePeOposHWrUTZSDU0wIUSgVecqQakUOc5ViXZH+Of3vkBiWZAHEbkB7rB6F+n9rPMyHFNUbI4C9O
+LMGASdsXRdUd/H1WNnC8utSuQK+qs91NpXdmHk92LxSJWm2+lKFV8rVFzWT6JijJ6HgQm6ltrW/
NuIhyMAPG0lrVLVwTd+rvgEekGkBXRf4MhmlpyRzjGwHBN2FRu+m8Q3kny5dOmTdpuew+JR7Uwsx
CWlsBAZSIcIcUjjTvWHpszIZ5LxBQxpt1wuINDqxnb4YSutrnKzakqD8yohcyNgJPO088oOPhGZa
CvskHcswm0Aq6OTi2HR+R2P+rpq49iB4Kn+V7XNBpbNYf9qwCoDnFNSeU00FHxN7dViky2ZcU5a1
T5dY4NwDqbpDXnJOnYmWPfeWz4CqMABwyGg06CFzylZznv0t6tOJYGdQsfuvqVRzU1HYuK/bgKfF
9+hUUwl3gup98Rzao1zuVuwBHwvTqovOT8HmzpfGGgI25y8hy6Jhj1eaDlqhDad70yEy+MXLdgPo
BmUGRWTTxMGA0ZAS1LNVKrCnsXDHI2sLTEj7ovIex846x5UK9V2WQPaS+7J9e91MYqCQdyvwV77K
bARt7UV38mKh/27iEo2xemEcn1PqtywZv6JF4FJztTLLOinMikynGuFyI5AVXUksjrAosqICmPQO
/+497Z8FvsWyMXrqDWRK973dZpOIEu2Pbz8eOlnqD55hG0EsQjm10Z56zh+J/lz+5ICI4I1q1rXY
spGRntrKgliSFvHiMx8TSXcsp6NY4RK7KxFqeSjE/fWz6XH30rEnqQsWm00pLV08OwZdhNlCUkMX
cRf9JSu/Uaa9QUwNbQp31z+U7RDc9Yz0gShMn1mwLRdNHpCy5VYl7EU5Sf6Wbc6GTXVJ7A/19D6R
Zr/pA4r3fJlgD9bd3094GZLKFk8nKJCLSMQbqbnwvJbCPUImYy7i6+OnALt7rWBVJX8l3J/t/jaN
DVjWtxw7IeZ42CVNhRWp1aKD/BUdjxqkCTTyRjmMLB4iTYDY4qDI8iDtlsMLNOXbbUjTBfl5FRDf
JmxOTeVytecJz9CR95/PkAaLD97t0Tm5JxinP6eh945fd0xloc1OEEC3x8qvS+ikFJc2h3N7oKwc
I9cTTp+PAi1wbhQOVUjp+Q6/0L119eDi5I6WGVIse/WFBBIDN9GF79/LjDvJx7gbF6CH/HA/Yrni
yWKU7rSS+4L2K7ENFatqP8pjySJPZVcfs2Q61HyXWH19OSEq5oT4Ij7NiLK4Zm49pLO7D9eIeHLd
CXBMEgAfGRMrEe8wwDvkVsKxcWCW/sb7oT/Orpoicg19zoGr+B5LsE0OXYfESY3n43Xm6T5i7oQ6
+eciJ7np5MpBLCjAvjkdyeNRJba3QA5pO/BJb4xxjXsxrmL7/FRE0KEqHIakCZ2Xq/4d0DCK5Hfr
JUBhSb9VuKNEG8sGK7zpc6yScQMYcR1a9NEql/i+N8jqHdMOetzs9i7i9wTpNJbYc1xG83/s8z9k
9NWE3a3J/m5f8EYkLJqI+LljxDc5ALLe9gn5XS494AV+VVbqeOpcMOPQCA5D8Wh43jM7gd0KdOq0
O+sGEyOh6njjE8VYdRGheDBehW4ocpQQutbDGkbrijDI34jPF7hd9VzvGRsHIU9ALvcK0Tr8QZOY
4UddRCcLx2G7A4zZtn1mq0CBzhmdIOHi6Ab7oUVjr8FfmXxClmXRzNvVlTSlIad2KZicBSBKHNEC
DE0ZrI/VrwqnW3EkOiZEI7ArWgEI4hGXZ1Qr519xjH8x23IYaBCiCnCdxbkvgtNP6xC64aVIUuAF
evJDIJHTK7CxskwbpjI/aMAM/PsL0I2sJOWUmIFH6EMe4d+UJDb2HXrx3oE+7PAKbKtKvOhAYNCA
SdgYD4NMFQl9JmwJghmSHKAIuVzomApgv0ycExdBgg+wUndmD1EZMLBhdhz1GXrYkzKoPZj33j3C
CHbJhXxx4M53eQgP0XafFP54bSXN+I6v6mFLnIXDXeOlSq51auyR7Q6mzSbxH5ARAwjaj0QWIH79
U7vzREX+LrFdIAsh0EeLNrq/RujC43GxKHcGCeXVKaq4D1cERTCG0q2wTcSOZlzzS9k51jIGni7t
t+ib2XoOqTGMaJyw5wTuCQxIM48YUpaO8cEhFOXLlU6/v4cJG6p0q1ikkPGO039n0D+QP9h76A17
WIawiodTUdLwQAp2N2RpLHhGOueFW+nPPjtjBwT3T+g1nmRecx6AMvb9vhKo34YH+KB4rQdXTrq9
DYtCVklkNdx6X6FK0YGsqD6iSlMiX3TBS2LVRC9zKM6NGAz8rOY6papMX11XMN1tKL3jnEO+CzPd
6PISB08EcNyqxDvKwVhzA/hbU8/Fak4Iv7srUWpGrbm44oW0JHvuA5MNvNs9V/vv2g94WDDtS+R0
QACkm86PymunZL1Nh4uZTZRkzuw6b286YXo3Av/CJ/Fbdfye0J1VXYJhEUBM+sgh2RJhTG9uXrQy
fV6z4dtNMIOi+iPd2ehgVJ5Y9B7DjJ9wfPYLfwFycgYtyV/HrTpOf9cv1MuEBHK0uGS7rHJ/A7/5
1FjaMmGMo1ZIehOhC6lp6irQotVRdlhI9vC2uIjVRVwSfU5gMbEXe6t8iggm5dwylGuXe5cX/Pxd
2OvEPLLb4h+UrHd+mM+k5v/6vQpARNZrTkZWAkrivP5MR5n/qo9LCGV9Ck9SLzo3dlOee2OKiG09
JON9cZQHpdVrn9r7mioGXD1fiLmg89nI/TbkIdYusIXCfZDRSCUIh3X8SB7rKZq5oic9ePZyaWxb
x3hdBSmFvSEXKroBm6dboEmttFFMACKnbuHgdKdaOFFG7ctVp+J54TzeqPP4d6J9wUAf4b8sfdKB
m87ofSv9MptBvpbyhmeVWzCzKGJ2x+b2qZNcsUsnfeohXWz4m1jTc1gvEVh6iADi1In7QilUjT6t
9Oyotd8GJc1r/Z9gVGnphLJD0W68g0rf+fxIaMk2jCqc2FRN2dogmiEmpwZnzXTAhJaGZy9Afdy1
Wr5+rh+2FpIeIZ14q4pyOq4vOkDXM3wJS6RWgg8VdkCfv2pUu7+gBTOQjJ6pPtFB0kqok7NH7Tdz
K+v/1oepPmXaMvsL3IjgG/7H163g48DHApLjqagU+edgoR7dFyFTAqQxe6x48nxjVm8sUd3w0Xvh
fnxLDcoRW86q+t9aohIs5U+LJTnLvJ9D+59wNd/Y2AWWxAk+sIxJb1GmxEY41TleitD5Da+Io/zc
IHL4pILqfjuKQ+PRkBTDtvaEAq6I1eUGN+NQBq8IgMFlwaNKIZMv196Am6EYTlFzFcQeHv5YX6IC
BcVaMQ94U0ZluZoyfRI4QEhc/TWVKKrBi9qI/6LOxeQJfNM2anejIWoSmWKRZhTzsYHwidy5P/wg
Qa9/wBuqhYWmmnpyiPRVsYTQoELWre0/my3QDvywsrsgmI1wurN6HOwBHy5zeqwCCNBskyCUf62T
NjNyuWUzcDvPu8GXqU5e9S7z2lLXClzCohv6b8VSF2SzlSn9awQcIF2/4TVGmbPHyMLx0rxEtSkn
3dqYkrhCys9Msa7yfMuY6DsTfj7IbjfDUIjhrnyJu7v6aPuDWWwzS4L95a+WOYXP6QX09q4ylmAj
XIkOcCH0vQx9LzuFo5j/kMWFg/9YwbC7IAbho1/TEoksAUuKrqLTW1oVWsLzy3iQNZ7vSU+hmxCy
/POjTEJSYOJHJvQqfjX7+lcQvv9lJOIP827xaxGXIxh4+YeqeciyeYQci97MUUs/kl9ZSE10za5M
Qa01dWHY/jCL9scZOwD25ylw4yeGjYMcFbThEr2qb4eYxay6UVwFewpspSYDR/J7TvvhroxRvYzx
yoMck12cvDPKotAUviKc/iIBPT04zVDbVFVYssSErf5Da6M/WWMQtc4gQggwZ26TiZ2ZTXuIjo9V
CwkqdoZYSWfjL5U3P2U9vao2puSfoqVUeuLAoSHNf0bpisNJoQbxg45TiVwT7Ht4PDUqtvBcvJ6J
Bexnq2B4KkuZxc82MED8NLL9ejO047zAAEae3CIRjjCf93aaCBgiNwX3yr/UDyBEnr2U0QeIv5kF
ASFpM3OPEapRkjOadziDjrKHi77Qiwd4pC/4L6+kZ3MSOh5R5fsdzGc4zTd/Ep8t/yRVoeXua7mx
XEAXWa5xKHsXbWvh/cZJGOgzUSbEcZqKLDzlr9yg993plMkD5WfYemRaH5ilnacGmwKf1NaYl5rt
3lAqbozOxw//x2znFQTWU1Ur837SRBva7LAYYcSODqKw9S6tVLQ9Hy2gkTS+ON8RXojKIgHpLklE
KyddlwANeQxNPjfq78sf+0opkeJQlB94SeufsIuKaFHhCIbJt5gsDMwOf2Sf2dkzC95lSfANvJWj
JwTmRYQQ5BRGQjwbRJdA6JNzXIAj/GZDeEZVDwjZ8938Xt2lKHWl1D8HQQZWkE3wZA8IsuybU05u
m8ODpmHZ/uE0JWfOMpuF03h5Aqm4uoCPBqGutOwt0L5kfE5CKn7K+thkbq3Mz/cTSESMQB50/gji
KX2u4Wk8fRLIxFOXMZwRmzTjq5GpGiook6c/rgTqlRWAHQtO2XbtWioa7I5VNd0MyuUgI5S3H3h8
4I8tbgXEAjli77CsSqoktNzB1v1gRHTuZYgT+BbARIHfpjSiWwx+mqDpjT/I67uFuBg2e8zVjA6N
eNBwDAAbQagQNlPfvdDoEZ0NfYDE3KBOH7haQvuC0P8cwQG6HopN9o305QCrPwmpj3hifzZ9qcn+
JIHFikOXgAehFfR7h6HCzKXVRv4uf11wjF7Qc4AHwqDqReOWF5BYLkjgB1ri0sETG48n9NG5boBh
SXtNnBl8prrJuhN13h5rTbQJnzheH+yDTndWIUSHhur3AOxxJWbqexDlDxMyZwQHP4C3mOujki2C
Paqp1iSHmS6IVaKKo66EFGLx2bBOPlvpzh7JL5QUgHZ1EAn5B3Yu57tvuhaDHB3KyA3k5Wes+JQa
9GYQ3clmOkYCAJuhHXue5vpUPH/f8IneHKbR1mItPnSbaGaI7ioUcvnmJAAx4AtByW+waFFk82OE
xdlSGWjoh94UyigNcc8RzFtL1SXrOzFevQA3bmpxZOI7z3Bm0UfNa/f4cCJ6reZ3/0GeCnduAe3j
ETsq0YahInrvbqJk3VlViWJQ362YqJSvexi2ef45/wmhsoYd/gTlJ6SBBSlByQr/JSscbCb47x7u
ooSDMvJXNbh5aDWAzNpIlYrwL6ptqdEcekvCNQa/fFfdLKKQgIxZFIxYNM+dS2ipLi4/b4IxnhTL
bZqTRmxRehqhlf1uFefKfH4kcNbw8ziRodZwAakKL/T/WzYWsFGX8t1q4FFVhi9fSGgiY02qgVJB
B2JqqhkEeXoDjQS3oVPsyiCoon/zyC/l+8MQg+ek0NwD5DcLytRL/m6GAzuTKpyjY9pIBBOvV+h+
uaQ8Dhf2lsudUkRyJ3VN6td1tR6t//JOuREo9BpPnJJ5UuikByI9F0zrUGWcyqiegyCCA2oLQIVm
5d6iDWAOx4eTCeRsuitpDxEPNcP/1tWqTWMvMPm2cSFS7o4NKyzlr7Oc7zuBqBFH46D+XtzyqOwt
IwIJKULhSwgp/d+YAs1xzEmvEDyu7ucveaw+xlLbj0mTxmI+Sbz3z9+V7yUg51SDitYKbFJpSyvz
e5NL+vMSTX8ZLNIFZSu+gmEQfDy6vxFqsiXx+fAMs3NG/ht2EaKxWd0snV0B37B+hXj4tZWixViV
t2VlxDPwDYiZ9hZNxJ9I241hAoFmbXh7YF6MK4LEEf17vHEwUMmqUD9J5T8avXl9rt8pVoDFzcDj
qAkQyUNu4atd/C99AXscwZNQkJ7QgKy7Utt+edmzPtoLiDrmx18IBTgwBNxBvVNDPxfKh5QZm9g5
bjBDSENiqjadaDh235S0CtTjj7LdpK89y9XQXpg4wop62vG0DRYRjJXKUSBJTLFEGZrM7DJsjLYG
vsuZcDLWs/lvI7em9SzZbZXWsNhAVRP49AS+CGdehAyLvG16ECuJzGH4JEESx2C5mOZeRGDm/WiI
1/K8C3sgWtvv3f2hzChLgDhGaZTzmXFVfLDzn+G52r+56AHiprcB0aFdRRwijv6G2Wd59f/GqPub
mkJLAMrRUhXTu7cvy+Hus67XjRwDv8IrmSIJn6k4L3SKoIJvRvl9sXG7+/6P4rFCgYcnMbUk0luW
8E1s6yUDztCR3jjyui2pxy5T76B/wJHSr8TbwvODaJ945ygF4NqHn8TS7RTqbhr+RzjmGATNtD6a
ueHh7jiFuonFF6XfwCiXtCBORIbDXrJsRe+1VEVHSPfBMKFaKYEm14tGBmS33idlDihIs024RKi8
xBmyLWd5msaNXDZFSNvd6ZrXqLeFKWpdHOTMoRvSMcBJA5a0CH7TOe82DtsPvOTqYaAugzssGZ6g
CIDOv/KME2rqJOAZJeYJJ25vqwQ3n4wdpv4ozDFxzEYIc+vG5vex3QpPceNhH4B8L4LPHDdn8L3l
J3IeoNa6kAO1RKaDUc5cEFDOsZAE9dMVp0ZqPE1U5lHa7N5cD8YXqXJAHRw4+a/C8EUqceTmeOku
FgqjjSKJ9IUvvYlY/pNNCUlqrFsd1gFhCx9p5fEx5PwIZlOUufjAsx8gce+Kzc0RE4UAsTD/G+JT
cpX3GCt1pVdyfB3fakeHYTVWCC4tQHRBTruS1P3dd7fPSwjpUeaUl5PhzEMSp1HwJHYnYvgFQguC
FtLKyCdY5USA+8wNGMFqFa/Q1XmNZyI6AC0py4cGPjwgjPHbFQ2iRdNL2nz349XV2SoRrVrzhI2o
KAaubCiFES3Xk4B6r0pfYGoo/yec1Em1iY7wzky1Fcl62lOM5NfZJFeEIFTrBRqZkG4H3fA5MC5J
wxcHYLcA87ZHf2QZxdBvirht0YkeGOx0YHY7ovoH/okxG+V5juRTYp6p2hWjmjLVMqoUXzQpOWno
Zl1/0Mxrk3NiazEo2QeqAnd+R0L5m1WHLiPTjiTHP3KQwvFE8SZ9t9kt7kc/tSftOPA6JGYqBjaM
mMQYerYbSBG44BNdsiHdwRt5ZlgD3cMPw3kKsLUOS4thIgbyym5VwaDSa4aMAmqH79AodA4n/BZx
P0o1WE6Hr6mkFRLot9kM/yZYvX1pJM8vFpVKXLNXu01qg1Bkhb7faKfhMHgmc4PDCHzFgW3+ZCS1
sugAtcKAeoFf13pSgue4yA21AiSV22EwW/pM+xKdO2kII0H3xcbml4VXxEUPv1+KDj8b+tL4XqLc
ebTH/0VRh9Qq2r8YpZx5IewzunoSGNS/j4Pm5AIPByruyv4BP2kAfhjFjmHXmns4TBNynWpnQRdE
bwNw4Nf3LMUzVy78ZUtq7ora2OaSZNYGMhFn38haBJ0gQ1f7pTlgL6bon3aQYGhWcDq9nYEK6yO5
TJMErZHrEagbNW+S8or2xJIX/FFhj+9hKiZzS68V6jTRUBdAxW3r0TYrteUe5yt3hQ0JPmORxYNB
P/mYO+7JWBO8KDpEqHrLfokx0ng4xyLN8Ht5T7SqpvPl5ehqZ1mYCkvZ0RxxP+EeUxg1W1TBvTgD
6bS6StUEZzs+33X+bM3WCvdKV8YrLJF2HBDIk7l3kLiRVoe0ULWGD2bwUTnSrCX1/xTfs5Z8QK4C
SomwWj0tIB13b+hkNKaDAMFzVsvabv5nhUtxuda4xkKw/pSMDzJRwvmq4r3GiZFCEYIvlRUdZr/P
iDSEpBpIGCRnCrhnP/npdCl3ud1EW0VdH33Qd5iuiT04E0538ARUbOEN0sw3S5aJ8cu+cJJ4cd0i
k5ndczCnPaYWU1w5KRu0U947ml8h3CeLvYakQFQLrlQUD7elhw5/zOAhnqZ1PxNKwG4J4cHddT4i
arqimj0jFEMEul6TPTGefQl5VVMg4P6+AdQGU6YnQD+MSCfaAJmz620Qv5HC+m3+TYn0zecwbQqk
mInRXNeS8og0DG1frOlHJ96Yp239de0+AsBWWbH3oY2PaZYDol/GEJGLp9z3hBwp4pQDqPyMkpNe
G9ebrm77hPNFsDxgFSytHBg5XxjSX60KMsDA5m/foMllsHBx5ILYn+xtu5DGkrW9zIP6NMXBYuPn
M8GY4RdK6WROfpqcEZkDyfc9soClWsop+10pJ03RXdaVZs9ymBmPqfnpAuup8Qc134byETEoU1pW
J4c6ryLsFQEMEbcoGQGHMXrmkzqzzhCt6IBGCtdJY8CTeo/0GQ54MwKO3T42WwBK7GWS9YtJm928
AbmBXZTkCWOFFzs9eM+3GDGeUB2HpQalvB0w18QiHwwgm3Ire6JbGs9PIehJR5iU54BvO3RbjGwt
sOlyaYOfHyTDaJFw3j2WKURwizOhCMkk+B50g+H4mFWAKgUHBZeZQJQSs2WIsHyB7yBvvtexIkV6
dvfwj6ehiIZTW5PJJQffLT+VhMUjSb8+rGLG0YigyDQ0VgYyDP9qlXUJbm6nzH7Xnciu6tTf/sip
4frsBQ65XRMVoA640diHD18S4x0ukjZq3qc0WB1EcmUDgMJ90MGE/Y+zplPJjqS52FIKCHbcrAL7
Apenm1vBeYs6INRWUtQa022QaTBjyJYGRWf4uzsZUfD/sZ6xd4g5Zf7N7GLHOI68wPRQRjRzdWJA
7gbQ39VDz5iBkkiC6dl8KZEpJDz1uT/NGdiZFjRaNKGQGghtSkRsDuJ1wog1GvHWLtxEH4H6o4ss
4c3HWAbR3/MWOj9+m8t0+4tGAjVNscOpJWx7m6WD1kifeTxd1tuLUJHOj5Q/QqYAH/p/3gsvKolf
ctKKEzu92uon+LhwSDd93QzqXUCYRBowQSDYmgOGhWRz9B7UECefXedq1SpION9ic7uv9iPVqOFR
gOyb0SRNGIo8ZDlO5bVxvi82qFxqWuwTFSAeeqynQaUoXk4cpzpX3MV/pm2a/d8aoTrLqpEsCuGn
ZCPcqJp/pnc7X+dq+CQFAWddW50Oh+i71NNSYrpmc4WJn88CfMrmik3U0nbblZoz2czOJLGOyY3/
EhQh54I1BV6GEeIRL7n2Nx+tuRHULXpAjcQvk29GXl5suhASWbPcscL+W8iqFnRWpJxKYC2pO7wv
IbEOys/XK0i95xT2/jdTlUGgGEJ9bb+J8kxX5MVXuRWvsCzlu2+MSnuEIOMSJ9+PFZwDPyXIU6Gn
BvSRnQfmnUUWm54Fq2NY8JpAFNI3EVVob2jZKySrRBkAPNzDM47PoF/HKb4zHjouS91UE0JW5C1r
pCkUpoCp/o8w2ZPb1SBCnscHqMsfQgFNSbizFAQ9qjLp5y5IJdHyucod2v5BjJhoV2h+5EbxiP/W
4Ky38zNuQEfuxVsWKeE3gB3pN8VV2y9PW7dNO5aQ26bTlpr9AnNRDECuDbPzEY+02T0vU9SlzRNk
PhQkmtUsvH70vPs7SJRBjE6onKuO9DYg+mbdjSCM42bqXFimtMlRfRNjJyRGmN5+LSdC8cEkY9IH
3OGW79v4ZGJOUQK+A/OFd8ClH2zGF0+7AChEsd5ooyi75L3KRVVo8xCYCRKR3cxxuIdf09RwujMW
VzEBV2zpdZvZOQZeunnVF8r7/Pe39ut0qbY4l9Kov8XnmtmmuDLH9WHkc7AocMw6A4XcMmzwubkd
/WJPN8ofPzA0qIoTHZVfKgOMve4yTiFJBb/6bP7XTI8wZX0DZqRG0kp/ku5XmeFpoUbBOz67Tzcx
uuXjOgsOvl0ATBNDfxNKdP3R66fadSWEYEGollWP/3JvEwb2sF3c0xYFNFgGgnLo+7SfNftJ8oCk
RHVTlOlU6lKks/VpZ9oYNO9iQef7U4W3KyFR+XOm5K8fhHoKrP1UKB1gA/zOv4Z7Hg0Z0OQaewjn
t831AzJIW9D4gl0h/bTX0WcMOZ20LfcrgK5HZsEqHGNhGa9/9O0UmBE5fhulgjiXtpu6wjI7rJ0d
dDnolWE0DDOUorx/QJfsPQp2ci76oMcNq0XR1ga6c4PobaNCrJqprMWyyL1HVvsqbiQtTkSSmnRq
TDwLQ9wjUntnBEy0SvyiLL+UjvL9RBuNJ1VlUywo3YlJ9Vv5PZOXxJfU5Oipta7WDbc5Cm7D1m6p
oidM+HqC+niHN3QNbLBb1ru6qQct7I9ufu4lGS8KsH/D64jcVUyc96gTzRbTTNzH/a0PLJwPCtSU
ih/mpR0sx86lvQp+7HVDxg03ZMtwOMSmyBYMdLws08vLBaNbZp35EJh6OH8f3cF3toJileSK1f8W
zCXP9q/dFNW59YXMXJAwA7aACxKq602Me4AzpCVT0B48kYurpr7TaS0nliuALXxpwwltbOfypzWg
LBIlo8lMZRxwMOiufUhIFQyn2tqjv1m4h21E0S2NV1kNot9QAhAIUjM9LUXdkpdwEY8hSM6J87TK
krrCr20iZ2MgcOm1nJVN8pmda7Dtkv7d6e1QidyYiuLvurbTucf4osBgZwZv4gAUl+gu+Azje/1X
O2hbfqYwiWETI1FviPcR4aBhwuGPn4xCtJXUB9zxNFAW9TgYQtVFofTuQ9KNJgD01uVcfbvhv3CC
JCnKBL0FaHVMyLvzRhcUiIbzVwLvo/7MjPNlJjFZtK9A4Y/4PKc7zARijV8edPu7yYqklraZ4T4R
Oj4xbcYk+dv2YUxJhPuRpxs5BOkf2QDqnzjG1T4vY1nLdpxQQtEmt4WNyHX3ATdWIaUu9JW/u8iq
cTl+LaaZvFay3wh81NZcrTnmQxrdjQ9kysrrmPIWevXnAYLM1yoBGgleV5IEdaFjm1XIOu/UxYPH
O6dW2VamhGUVdA6GHvq+SZS30u/vdtKb7H4Kn8slCarWUTqDpiw/HG7LECukMBfgawPDHkUehM91
gTtYLIpPrAAo0wwBAgs1fspa3BSVaB21AIs3oOXbs+BvZmFQFRDY7XzX1cCnlTXA+2x4M8LSj9nm
5pSJFvHs/zFJgut/PtIgVdmogCI03Yen6b9sH7XOONjysbuhi5/WrXH1F1sQkBpkuhVSxXdoe6qb
j3AYKlc+URXLabgRWYwArEzkWIuh30YtvC6D+IIRtUYTqPlccjH+JSS112YNbX6KuExR8plJdwKx
9cV9E4ix3EbsMO5O7dLVlAc8rCK8MLkp3DqGDN19R/jugXWmqNIkmsgTmolWpmW+wgx2xb6tJuhj
STUN1yNUXywB7ZL0evOJE0YoddPEjFzcCe+vl21XylB1kYme98fabXlMVcxbZ+VwqxE9zujDMArE
golQfOODjAHQqUpGNzHhb1S3aAamnCB+f8evwyJm4VtglXTs1q8nj1FW6Putmg9SZPmdQHColw3+
nDWdXkYPcfG4VISxfKSOEW+3QkafVSqAs/OhFYdweBIQf2x35S+CNnDEvPO75A5jzDjLgoikzi7n
IDTF5WcEOajW0eV+ejXtPfDKewOW9y+rgmOVNDhIJilLWPOmrOguX/h8KBeSi6vF0qd6c4L4pLOY
wWp5WngIowueEbz7pV9i4mLIFgCMVIBnnnqOn1nymzI1UqccAPm2rJ+a+hQSPi3hl1NvDYR+i4yb
y6I5THFjtkTC9/ZXaeVD6J4o7lBbCArsvBrCXeTxGvLu6kvZH9g0uo6+lccqx66LfxTz+y8LWvTu
YaYohLRN08GZRe7vOMMf4u/oN1SjrB08yE21/4YBQ4P1zO3AtDPYICicti5KLnS7Tis1WmQq4MyX
bepOikW2UkmFWP3aChpED3+hpSwXxNha30ifzVHOb4NK6tMOzMsM0akDeMliGmQVPr46Gt8E6Wjm
KVYlyrRzX6RyvMuhwxK4KJxw8S0QivuIxTugbGA1mUybsG/GrG8aBXta78Ms1M0ExjyVp6szrYSm
BixtCOCLX2emkQX0uJoKODhNWzKL+dFwkpalDWb3C/DHzmGDxjKJeN9G7kSh+6ov6yHMgXpfNiH/
1KBH0v8iqhzas2hYAZhs9T6wSkE63SCw+HIV3bfb5kISlQssN+7Gv68GeTaU374kmjtQogyHpf4m
Td1pO2Q1oUpecFJuq80h+fxJBGX9d0/h9acHCJkPxuT+SwXNOd99uyU2vePCbWFBqUxy5APHIAS0
iFIPevzUmELzYkFEIWzYxhhjeGC/2dLpxB/LQKOXwz4o/aljJL0YCs8Gm9nvyp0GSDcLPWydr+T2
5xbi4o23NHrb1sUp66BcZEFlm76p4tdqVsEVsTs5bFSEmbfRFhM9W4/MUnHTw2nWrxCe8anTGgnl
UJyz3o3Uqgc4vKkdxE1OD43F5MGRiW29m1FrYGr3LUfLYjW6vDaSCWM174dFuHiS8kf6PHuUOY2a
2o/QVmk5t82Lev8pv5JnOgRtaDkiMddvFakZjDvSpXEVhKHH7siNgEC9eWW4rOUZZoXFCzd6dV3N
Rdrga0OSl0ja9VAsiKXJhsWC4kp9LaevdNzfoDZdBbKrcoqapPRvWnjqrbZ2BgxAooM3kp2JrjqC
7Xr8gRL+2kZNqAqNWVLMZmGVuqC50SO3qiwzC9OH0Cz4RLbShOVolxU8KPgxGhxaMBa4heDyTjEE
2zJgKP1hjupO8SOOZtJJYj2E5vBPS8Z2X3+D4q5n0yZBUXnpdwVb6S+ghpNXRSgIy1kMU93b7jRe
mKUjIHQpCKhPpWJbTlXjSro6EAqcpDAZWorxJnQ/LqvMWGQBb643NNr6kCu6lIx0yC+18+uIMAu1
biUtvFzmIR/mQ1hDgoRAtq5R7seERU4QbvlRGAuZicsvDMwR9kk1OKRgmHuaY3aidmI42ikC7PN/
ocEwaJ30KsPBB8nreuNyXZob4aAL/pbVkrmRydObhE/QtCCMFjoq/b2vnF6b8Ne9R+dXJQ0w0uW7
PpzulaE6Cb9ombUKk/vXyzxGEMYmpOgbiivs0pEOskkoW17Pcl85+rULkVUTV14s6jjnrNSVOE77
w9fmHgp3qNF4BnI8+JTWWDRFoBBaXdROucYn/9BUfVDj7JO9DRqZRRI2hD4gkpbeWIwPmGjJlmDN
d9wUEb9rkBKOIFGGQvYXolU0yGIzT1pWtsUpCeeFssMb7T/cdBPCcqyP/roqVavxd1c6tYPNI9uL
F6BpgiPU9im4ZpFM25dAs8UgssDcoT2qfdzXV79p5SrnUpnoGGJnLK3UwQwbb6oFwKDfJCRs+6mP
3ciHp5hvpb1CM3giPI2cOHvh0qltpVm2zOcFuD7ZPGczW4bvy6nzzkMCX3I0NJYpxhljaWk82ED0
WnAAM/T2LPyaama3tVle5SpWI4H+lJQ80JvaYuCZcITCoVdDZ8+wjB5anoAEr2BfWfSOQblbr7Fa
x62tkd5KgesjPU2U+/CGyJBmfK+uvOAGfMrQTImg90+JnDb5mrUmqLRZpm4FhD59JB9TSsr5eH64
8Q9bdQIY24HP2TwrszJ44dU3jcpqpXomYpoK40thCEe5BfCpknzOe6k9IKj+4lxGqhi/zxYL1zFU
sorYQ1rsLMYZpoJOwVMnsjQvzog0yklxDb7fQPpy3R03UhRDBtofO4ESPMm4o3Biwfvnpg83cr2/
Y7P+G3NbQgRw9KX6GT9sgGefFIOD396URwBx+MBdXF2fwHlD3rCDmwOTph/aMXFbdT67pMFvOPlt
p418s5Vjp3thiza7oEIRRrp70MaD/RbTqgRFNdLhdxSwKdkLCRHGGVEmryg9Ubgp4o6ukBEgZQO+
zL/upwXxoMBTJC52SOb+c+avklj7fk/QqutwYcodaSDdhPLt5NEvhYTRgQIsM0XhB8mGiWB9LPsa
/naVMNZRFsBWHI0eX8sulssfBGGm1x2f2x31Cvgx7Xr3e7OYzAesTpMCYHtsSGRkKTyKKTgpT3/j
25MhnQT+TVxcapT/tg9ECBXupm9i89aeaT8MxP92bxxyHrKLFiEUeah7YE01jYmukgaQRVmgcl6X
3P1/XOE1Vl5sCW1gHIGYhaOcx869XcBKuJo9z58QJtcLJQXIaqpdET8GPTYo50V4mRFhXaA2r1jQ
9CLxM+gAIBDfKc/u3GfxDRMTXujUJtgsMfeV4lmOI0lrYWql+D25f3KZY/M7pvtBADl/xCJj/7XA
YkVCrp/+Sz/JsqLdkexG5eVCxikvIY81WzMhv/X8on6AGQFdNZoLeUpGIK/uDTAhpIupd5oTFC0k
dDiM30xKEgOEe5rWBLIOsllOucynqxQEwvWKJcOHzUgrx5ZCf7ILv4FxlfBdfTF6ivaW9XoHqSo5
kcmQMYJujirouEWbUZlR/J6tCOa6hyjfISpX9ofcUhcKMCgHxry98CwnnKR0/n8amx+/J5tWYCG5
sCG66A22ECLQk4B8gQpKd19baM2hxcfE00cOsrLRHoQUTkN/Sn2kHsCMfhP458qaodV9fNlu6MS2
YFLizGEbXJ1AyigSc6YYboMyXzv0ItSawM2803QJG4quFoLL2ZJ85Ez/j/bZy1OYH6nCemwL4u+W
JaHDU6p3XjIQ8WKxvR0ZcTk1LULsuc3QyAZf1wrFw+d2oUBVvIZkAtXcOclExGm2mmxs26VQLcyT
QG2AKTT32fOf2+VN5I/VxIrhrwkZnEsmBjf1jLG3LIxItaRuZM8FIGmfhaoGb5w8rkQ/Am+MeF30
QKwOdvXYI+O9y2B6qiUl5aMa0O8yqKRKbFzBYmB09/DCLDKwM3/1KK43YPbPrIuJYys12w6Tqm3m
3Mrd+dZ6jwcl8qiRdL4gIrCM8crxYiDJt3+LrSGPQdl2KcwE3JQNpCDqXusAb306/Gl1e4NmQ1RO
COI0xgZmluJyGTQWohW0t19dY73teLunVLHl5ucgqFqOmmoNSYLWcwl9nJcjvEBgDc+3hm2KrAS5
1/4pmkLg2lFt+/1ngN/EJZzjBpvsMb3Oi2IjyL0igVRtm1qPZpyyqjPTZifAR8RDa2wMwWqg0zuk
Ov6QjmLm1v778E+SwOxS8pK0yawcTWwTdD+A0FrXcGyPSYrJ8OWajV91D6mdrQEBWp7oFCy8zhtn
jh3qBedqZiTrhpY+l/qwD8h8zvMOCtBkpuruPK8fvfvhyJSUWjV2z22CgltH/Q/21ALuNYxpNd8Q
lGa9H7Qbf/KJnqxBXqHUfF4YIgwJQbe4odPykGAMiZXgUa5aCZbMEXh1o9BGDl0bNvXYj2oxfNuJ
uScu6lPd7DZhw17g5wtAHqpIo/dnQO3tabYplwIFjFdDNh7V90lw5xoHtrW9iBXHmQpxqJbM1xXB
VgxwZ17niJ68+PlxRgW6SO6HUUvn9bigba7QwE5ZWp8UtEiO6ZnKSRJlINPbmqe2FyYRTolV6jd5
dfyGqyRlqIEKspW7te8f2XAXpscUSPUyiclpvGqWx3GBqzlFdZlPBZt5aEwLkf15XzQWUvPZPubC
rD4Mjas78xH9KiHZKms/j001vXVxRKb9eDps2+GOFtPfubno//WbZ7597kr+RPEBYTWCcVku3gkt
+bhTBpg9AkwFc4MfXvp5Kl6mddRRcK0aAVD95iMBMuv+5BNz9ImWUG71lqjj+Fj8ae9S3WOo/V4k
QbxQR0USF/SLG2Fab8TzJWuFT0it1wGdiJc7Wcpg45n+iEe7IXZBSCeIrkLe9dmmbFMG0XJIW98P
SeTZtAz3VY+qYYPKhzg49yWUe0W3zwVo8gekSWh2lCr56yPYuDKYoPzFxfnOnIZ1po/le6CdKS6p
CDC5lbQpH4PLL4TPvfBYD+eRX5udlyogYnGkRTExmQZ3WQo8ezoTDFYIdJbHVOWHxijyNrSI0dtU
g3ZFFlD4Om/yVcjDa9x5yh3tHVE9F3fWbn2zLWp6tzpaFNC9W2brHJAyYYg1kmWs/fyx85kdvlob
u7s0fxaSG/8pv6ftxsDVOa2UtgASPc7cOWZMqldvTcFaFAE5bHuVUT1eYbkTbfyusUHaTWnni0LW
U0xVUuzn7KKBkTlgylce1Mta7K1s5jIRcpIKEUECuqD+UlGHh9j7XMdrLfSfmf847tMyNpMUu8Br
lntFXQVH5Z5mkOe1WRZn696LBgUvLGlsBardQBYpFB+frUUXYsyYUdsRlxs5sj4yWmEavIIms8yV
LVI97CGCDGbDNSJKIsyb6YzpHVtrUogJ0C/5Fo3tIrFq1zJKIHnvx/Spre0l5IEbDxwlATsp9mUM
QkgC+B0481PTRvJIMgdqelz8ZeGMLrl8ZWsOCnVb8x5c0etyv1hpFu+x1OgeLZSLfZckV9+5tMoX
bIcrgBOWM4QnTOm7NLep4+ai99/HBJSNIjVLJmkC023RGYxAUhrHW4ay+4RRSYnKZI930J4IrfBn
ivyOqqAzqmt6WL4M+yPQIImhjCYJ7S195/pxDPgnN+vvnrDyDioiwJY5aB4LUYdory7BiCj4X1ts
qYtLzGtuHhR9m9mu7HlILzdcVNpLPhvrwrmWq9cRpRvbm6cVPTZ33jEhAw53hvD0sIFVNs/8tBFl
FkU9yUZOJzeaf0HTSofgBCh40YI19UOxr+L5PU1xeAcGXL1qm+4gGY2Ik3M/ttcA+V+WQ69OXZJ6
uilHS4n+0qX2JE8puWY1XBArId+XyEJbFNa2GgVLm6tzLGJmGIaFF3BcyrU/tu87UIB52Q8ZwBkc
mjAQB7oCeoHd2ERx064PMiHqhOyVEwdPc8vaAglZ8/rpQ6SsZ/7fWtQcnNp8O24PIWA2GqdBRPph
QZaKo2dOnGzw41488abBAF6bkh3jnm1XsEN7BNVFTW5Od4ls84xpr9/BW9vXORsXNXI7VM6Uw/8e
BizFFNUSMhyHiof/aO4mrP3hvkLkD/peWsOwQSTcoPI+AsZOxJBpWelyAPAPhdv7SgjXb+BcjYHe
jGAnF6YtwiG0Kg0k+IF6JqgMU5mlY7emJkjMC4UVsQbYbz3CY5PXF/XKvVXF2sFRVFQLhd15XgRz
ceRX8sCGBuw58B99AnKJciBVEglD3wjOxsb+2WcpwAODlmB6PgVW+dpV//GGOXttpPcAoximQvuh
TXT2ZQwTOpUklQgGsATGsMgQ+Cr7vPiIOUIbL4Kor7N2jF8C7JZFhd4MESvt3TY/KU6H4W8jWKjY
SrRWcG2FYHnh8eEFJt+39PW+98GpsJmpibdz1c5S8JW8t7br4VgxTG8nfoqZeCmdXPg138rRLF1B
i7PY5YbsgmbAhqbnK1GQvBubF56CqqunKb63IXZvMrexxJgLYoa6EAmKCqz0JxnzjSK5mDWqnLco
jPCF/nOOtvbX/hSpU2UDW8QcLHYMp2kl9hd7OmaplWXAkeLrbvEyvBlFE7s7zy+G/y3n2a/aNGPN
Wl1I8tyKhcBnMRhM/8Vz3UrzSU97cA8buC3YtE2Y9NUTUKu3xRWkCUV1nJEF/OYIrqB3NbuKi9gV
2qq+Ab6CtaLygnRVu+H+LeDSpfRazwgjoRkSdhvIxY54GKJRKbLHxcsHVyd+UJSiPIt6N2tKXT3T
vhogijl6L9RNtO4fQUm0my/fLikl6S6FzzcqA+Nf5kzN3zWnAqYr/X7WPrpmbwKUuktCTDC1WuV6
yKIFDadjn0riYNtM5w1U6zQEViZtxQdx3LjE+MYhYmqMnXYj6YfNqA7FolXrVuItnLRONuu6OBYT
njnndH5RrVwwN29dFw6NFLlPLfQNSwWMYNamJ0xJSJNA6XIQ8HNdqnoVPYZoblr+1vvcs/gYmEuL
7j7Iv2qrDOm4f09ZIjrpLT1yJtrz6gQbri8OosCaP/lzkRjC1t2P2ehOZ0hNn83yj3SC4YAVlYGa
0WNfXgLG9Dl11xEo1MQftzZZybrJbk/qL8zgceNadp6yvMCvvkBcESLguLs7NcPnHC021GITdE/a
K+yQb+QdKR+OTIRbxtdFM8Q970jRyEaSg4zdC0A/lMVWlYumizEVDQviK9CsjNz9AjfjFB34n8o/
/NC2s1/EgZiPtQ+cbIl6q7NV+yGlF9LBTmxnNduEhkBsJb6G/CEdN70G9L3YwecSx/QA3a3n4vvH
NjDdx3ZlbC+PIta/KBHr91ftbbGZ66ZoX3a+e2hEbtwJixKXiueNLn1kJ7XayjQNMFkmXGyXSbIb
6erjomAwbAX4rO9GbP21qumAfP6gS4y/nWW8krcKHwTi+nDz4wvHkihCPOE+pC4XHo07jZdC6rLZ
9ioFFVZXbnEklMaPDOZzQWVNNINxwkRhSEqlz3GLqYG+xrzVfqFd5DEsL5jJetlaBc23e9WJfff+
Rr2MblhcGdHkhdbm6rgZ3Vo3eJBpNIs/lXNoLuJKOzSYOEHSwL9K28qyaS3dWb3iV+wZeeXwE6Gu
V0BEDBPQK1MZbn/B8jsvUyBlKpFIeBcribK5+l8bEy7vHkulv9qxKvcfqfDBZWXiH+upRotxT9lp
KEhNQih51GyPrhLLYF26Xc5NA7G5ZZ5sfrftMBUal05x3RdhbSw9RgJNn9Cfc9z6gSRhji2r/QtG
+pqGOOwNqzgm6T9ftoGjLluIlTiKrszg1dQ9sn8sbaGV3FkayGNHLjuM4aV6pJ1JQU97ZvkaXGrk
XGeyCWnfYOZHUg6t5Je0MmjHCUzt2gP8gc2gecrwAQUw7zprf47e4XKhpfnj0BezNVPUOCmUgFZc
KuYBlrq+28EZ00PMjd2wBHInEoZtwsvGf4pX0N9X19W/r/Uop3vAHkMb/x8y583VSbK2nr4psdgj
Kx/YUqMOxUYWq312Ge8+c+I726fkkcsXN//M8746x/tg9Tuvz+2qOVtDJqpLuE+Cj3B3HFi5APiF
2ZcM1Pi1N0sBmSsA/iF873pxaUsXHb6x9Qy984OZrElHga0m+bKJswEQz742Fclrih60QMFYxh2Z
BKwbGO6K9PYU671esJ7sL6xX8QF1XnuwF7bBVYpjdb87fAQekeM0ndd4d+fr75iv0JrhPU0QHv5r
P+C6vPEHvWJjJYBfaC8Dme1ROLtGAQaD9J/nqpgiGCrti5gusvcD7TWUzWqui9UqZ3Ug60X40kut
Qr80iA+NbBCiwLCGTLm/4+MW5JY+cK5TXR0s0D2vMsQgUKAO4T+V8BOhLi6U+oNoorYm3Ztb4UJM
JhR1VIpJgKChLwk9ey1oYE/J+Tb04g0kd1mTp8JL6d7kiydoHR3tW5W+dtTWfzvBXLjlIfyyW0M7
C+lRCneBWOqWjWFR2V3NVDwySpqNj/39Y3jemMKmpuIZSEoPVsnWt3AWnVhbEsQsfGGdqw+WHjae
w3cV9U0FOTRxs1ycWcvZFLZ/TCdGZMePqHQH8gh8jtPAv9ysat3YUCH8h1h3AKW8kjn/tZVhdIxO
6Mu6UvbYMFuY7AmN4o72a+S0S6RWQH8sSTZER1+m4WVSmHxvMslh3wCzzkqy4bvLXhMdHiibtVU0
FvQpSnc3AWIIsD4QM0h//jkuX7j1oiCTqfopEc5ov+D4L3DZkRcvNCaTyXPfmg3wdQM+i+dWrmg3
SdRjVYeSas3Wbw5Ik/3CXsc9ky+dJ0ow03Vnif5zzLy1lcPvvOpwjCXJ7TY9ac2NMZ8znPMJ9g7h
DcaCPXdD5VawkppZRtcBs7syya+bJwjBwf0G0Sj2oROovwTJMmqJSm9SfyPDFQGd0al5UQU4tuCz
mcSnJYeHYb1HEILtlSZImHowGSUO/IM4ICDaXvsfC6mHhGLBj2nqdsHNJrJzCv3aeOzRGyPmDI3f
qCMoAHY4CJo3Z0txSPOu/XLv4YopK+GLP44+kN4PNI9fkm4j3qOkGInMleoAD/Qz/IfUS6JjWmR+
72aORXvhwfzRIZV6RloCMLWLy45J0DRStjEg62zWFShUJEQqDMnMMAJSYjSTZC6y/L7GcAbzZSQv
3BOAMVShaiOSPnIinTiD4DU4upMIcp+RcFeJMug2UA+OBNggRsuqog/hQn0ii6O4jdRQOOx2Ffi5
fjiSI5YtUrzS636MO5VLqPf/Rg7veb7y3dI5rgB1hvpkGphdivcQM4bF/U4kDtdZvLW+FkQhJs71
jdrM0mUv1ypiOJDmV3ubQuB1nUWa5fEDSmwOZ8ME46ABDGxPtZlFem3gonhv3JQ9n/aFB2oVXpLb
9p7Q/cLL8nMHPSoJHZ/QLRlCJnBtAiVIrDX7fklvf3C5AchASNzcQqb8qRL6rJkThFgCpr2A7VXD
GUaXIPKObMaTciCDCcms07QKQd6I7QVA6CK8n02xVo6pbQt+nhB+ZA44tQSxYyQeGiJnELvDess/
2Hrr0soIXZva1lOEzwR4ErGqDZR75cn/0liDa9jMvbvANs/MoLrBdRYnMof04QmmdZf3irYPlNEs
ek/EXVT31BSgA9GEmkT7ezUrdzbJai5WZoldgpaxnO8ejX8f240CUSHvfmizPNBtSDaJfsEPupJ6
NfyNjRPUX3BcUeOtFDI1TVb2SRNIP20LkvMYbtDaaJ3GGG8ArxBb3tSBsC4q3wc6cZNB2VhLPO0W
qG4d3Rt+lGcglIq9k3CNGTrz1rIFfVJKIeYUS4owKp01jSsDv11ALUUaffdH9g451zbwlBwRdJ1n
qnEJzD6+4/tMtw+5sIozu3MdCV7jFsh6ItfaRY3TewtASLgmzFQj9m3FMh9wQu7pYKNOMQfiMC4G
jFTUcNVukfzsefK4rQ29/eTYxx5ij94sDhkrsYDMRr6Uk92jXet6DzCTuBZNOodX82Wy2y8p2/3E
PZfI8N+83f/1UUg5p+nES0AeWQGD4RP3OrxsC3DXsLHT80ULcZjkpb1UIrX7FfPRudQ1f+1VPTgN
k4QxHUQ3q9Xw/KVe77mHHZR3L9fwGt7iyBrdF6WP33xq9mWXxgc4VrEr72PuqEN8T6habFD1Lby0
KmKkmeutOWpvUERxS6ezRxW6brIyd7/tEHXtXG8c6hN5XxpomRujHtwOPKl5esJOGB5iYs0DByaC
cjLEtNY6fgAjW4IhBxGxIZLxdVaSuJLXnFe1mQqShhMWzAY8H7GsaPJwrbaP6VQZhIPngmOk3Ibo
xONB7xj+WWG1kh+E7VpijgEzaMyczUHjbHIuAWaS7l7pZVOMoF9p9e8UDk2WJm1ME4+pGDHLSIkk
iLlXjzJxDZCtsCPsHf9w1OE3L+DM8OzEn8L0PNcb4uH/gpZJO1+Ngmt9sTcRB9lfX5EEi2/AfA41
5w6rZY7nJmBRq9JfKAo/mXjCiGASoQtpu1JVBFaq5ccRvUc79nMM8YfXgm270aroztdXrGoKrWWT
xnVXoLzOa6q8UvnolbOB5tHKqT69P1VGWlj5D+UkYUp/4w38cUtX0cZQsWFkSQXcREgfbtpqQ+FT
ZIlFTmQpUZqGmNo8I0xSXSMb5QEb/hkqgxJ1Fkc9mWoKWuTebmgZefzy/HNSayMGAysWg0H/SObo
tQzjFrFClDHbM5SEsj8PctEHFnPjAHukZM4IxtdOxwSv43JjwDGcoxTspde6+MjfFZe/rDjYsqdT
uGVKCnky85Z2qociLZU6mjadisSEDjawbwmLsqXDsDfxguV2FJkBTV+zIl0haDz62pmLQAu4i7zv
/+D0H87srD3OHzv7DxhAt4/rZNdBYBQdoY1GEr3FVnb4L8pl/wwsdbn2Vw6q78wVjJ/Wnp7kNvnP
uwYWK7MkYtygOpde85RROpHtO20xUbzj90yjjC/Ri6PdRwAbEbB6YfPbQkbhmEA1NuI/5IQlE5IV
0EG29WB35PNhS6n+suziH6pxJh7W67AsoIonTN3eN5X+nWhyHGpHhuW+J8SBvzI3Uck7FLFCeb4X
KQXZxc7gB5M9yo0QyVuhaw9teAu3uvICe+3AIRUZgZG9+KcrIIy0b0XL83BUioHPRvHdDUf0e9CX
4wHXno+CeyBkeYMJSgoO25DNdYWENRS5GP4r62rqIukZLVsnpMd71Eky4Au/ID1Ag8MxnYBEzcLm
CygzAYRWPlDe8dbMuRU6+m2aibroPo/Uxyu2fdy9wFGzCTCrBki4yaGbnTo0ob5+7+0JH2JD1vzk
rsDrzX7Uf9SFqmaZYYWhS7Hs7HPdzh6Roa/QI/3ItMBLLzdqJ7VmJHfixUZ+HND/j9UTLb2lEHCV
/wRjh2A6AKOBULpsovxKNP8uQFm/MtstwxyQ71DeCuGXYalzMUVEJyBeicR398XR68/lSyQHe+Fo
2I6euefgk4r8ZfnkKyuq1fiTWxBOm9cOq5XP+HQHBVYsNuFbAK74PhllUk3hACfgp+zlsINTadyw
EiVh+Zroh4b0SQWfMKr0g51eK8goAC0/uImXn+ikv3UtlLYxEZDx0DYunPK7ixWjgWQYg+E6UL3j
v8IoCfZ5PfKEVgxl8N5p4Lri5JpvJ1fkYKQ8j4p+Sb8XmvdWYMaqWQCWfCtoo6Q32hg6GK9fa6dV
PXEaqNkwSXWnzCWGxb1afuf7cNfYiLNn43MnA47SToja31ACgOXPjwoMsgRQuxJBuIr4HhlFK3Ie
iRIzqEZMKTKUZXSYEZ676SlJD2QZ5aRku28mCMCPF1wKUpZgEpupNPhFKkKM8ZJZrhTsY4ByRXhF
Nu9F4RF6RbulzjRi3kHFLugdn6TH/owmAG4zjZ3go5iQL73rK+4osNutbrzhb9CHWW/y/bIKXEDM
vhq2NX4mQII3ZD3AXpVgVHYkjxVzEQWlEPXZAnXytdwlTlX6x6uvp3RnL+NhhhqhQCLbjPDn4ljZ
oL1wYIoXaW4U5vtH5/Bz4KxyQGX1qdM9Mg2h2Uu+pZcCs/9dwkv+EPJjxjx4ftSNuC0p5lklNRBs
jwLkuSGmGIVCAKLqPSK5mB8URZFekO762Cp4cQ0urVuutD+jhNd5xKdaqboVb0Pkd7Lf8gy/Eb2K
tPfw44En105sJJa6wW7LlMN7f1HVbIzXzzVl0fQdhWAvSy3dGL/j2xmKVPbLwe7BO7XJ9V1AJvfp
7x6ralP7HqEkxauxFbqsxtf2WLFQpklpE1XxZox2g47nrlIoEtZMdK2tkjZzZ0eyJK2d+tGoLy/z
obvJkl7TuzXYHrDszL/6mHzQgeX1gtOD5/mvQxl/J4xOL8JDsa0kN+K3UD7neNM1LnxQAlgt3qxy
n+7cjNSurpfjCIHb6MBa9/nh1tWL4onzCMamVdcKcSZnaO6Qx+XNiTo0kZu6ZI0vkmGC74Li6Juq
yqM6ogAJXP536NQhZaw9cDqrRdpk7UEIlghtaX8Et+YESJy0IpMshXU6aH2cCda9fGPenllclSE+
K7i6q0s9x2CVzxFx+t9vEJ7VEKs3JWDQJp2LlsrxK2s+n6CkUIbxOd+TojiiUk0PnFhqF2n9X7vZ
4Dmnw/y5CQkgmB2EUXVV8Irhd3DhWWGfOcvb2f2pxmMZNlhyuYPxrYsgWTsNqTI0ZLNKclJFYIxD
CsnpMKyqphwt2psY7vXc58nfLcQnba9oUOLHrqHrPza1ukPzE1llDaQy0TsEjORBOGIFOqItTkt/
eWvxrXcjXU2rg6QodL099yHUnL2KVdZItpkNCIGF+90/61inxs3CNfacOv9YQ5em1fll+Euyfcdw
EYUy6fHjkW3fO5tW4UENFRLEi/Jx7dXOtamODG3JrBLACZIb3noT0IOLb3erRMTvxqIqhZ12oRE2
YESK4xHoCnEkJRYkqRcHUr22oGNM/SY7Z+B7CanRMjcydKr5EMwFmrpCHYmMbtYOci84ALG8Vd9a
d2etLjdm7w6oxOHusUkfQwWARJgoLqaZT60Zse0vgzQ1psbD7i88Vm0gK3mvjuNitqJwOyHl2A/C
5RoV1WXYUtiMAffbPi0x+0CrfbU/ZWZoZeqORwIdRtR2sRDgnA7lrd8Izy1rJt01Fqr3dIUCmR76
5u5MYKwZc7utFdhlyuRem95Dmab15VHyh8NkKJeVsHq9kXoalRH1Y7r8OCcGTYUV4ob7rABKEmdz
oi+TeX/Ls9xPptcWOEQUTvsJZot7XYYlancNvzAH9eo8VBXdANOJ0j8ZxlAo+Mo9eVi5DRAEEu0J
hfQFdddRt7uU4jIUORa9eobIkkW6Bs7oeqp1lYDpqJfWkbBYI1p+o7KScOgBw6k4lJ+HF6F2pDkO
YpyS6higoRSDvmkmw2b7Y0UbyI25d8zOhmj5QL5V5TihSw9OvHt2IjanDT6g4CACmpJ4uHfjLROa
rahsDGMYHlH9wr9mGXFWBpggVZAiMJt/o/8WB8DIHNYhQ/kB2JMnSCtOBl2Oc8d/w+nCMTmZpDQZ
EOJg3wqifDkLPuYHnXQDscmeXlu2OjqctnUf8VL3WfvPN3SFHAdAR4VpTCewdepd9MBMGUDS6oJF
RLrr2Ae2b7K+BQEkwGM7UbYiLUG979cGncc+trCfZAHijvLWOQfp7CVbeq8bTp2XH312l46AjxtN
CX1gpDlZygTWsBTtnbXXmOBhZNpIp079lKPDrgS8QBpMwNUwDNQnLPexYkEm0/lUalqY/ac3xF2z
WoDSP/UA4F1cM+q6lPD+460pfVaFAFHJYCO9x1/38xX7fZ5ZBRavMaG26os/3MHkAkkXG968cNWF
lEU5SBOGRBZ+RYnxkdGsN5Ry1y4TFlh0QETPhm79BajKb7xlKrwz8k1hMjeFr27GoxYKbGVYLjlm
jvG8el7f8bLtEqA4nIoAcZuJL89ITkQ4BDruIgwkScysGd7zzOY6Jj03uRVs3f3ebLlCON2u9afE
OB66yzERcA63AQa48Nmcn/iMv42wfVfI10oM7O8shEVaeAMlXQnI7zlFl0PrqdZVJOVv85Z3EZN6
6m9Ys7NDEY/OKTikAw8OCOcBWmG1g1VOJPArKL/7Kfhg9ssS18Zxl1y+eXaP51bnuWqxkn1x89ei
Rx0pwlPoXj1bpqdlLwG6PkoVkCU598vJRfl7CI6QjZpvrXykKinRJLyDglpIP96KseU9zOh+xoBP
Qw04LOMQtzIDLNvYNUCxD7EFP6JpgPcGXqM+08FSv2NzXqIUop+VWmL+PKVsQypMsolH4UNyXiWu
SLLQCCPOcbCMux5f7XyLpk5DFF7vbPjo3uzG+XJLhT3zo0+vDi0yc3WMa5ZD0CVCvK+AgKdRAKU6
7HzbOkSGkfFLkNNDJkCLoWAK7vUQmdIZYdImSFc3LISCl/pu2rJJZltph4Q7iobqTjKVpQ8f7DWD
eWudJBekPIVYsEAc8BmHxAFIHnZVluEaze1Q2AD/BuDbMcdW9HOQL6H99eTu/XwF6qVFweQCu+Vt
Qiq+p3Er7JJ4+4S3yvzHpqIW4ufSqAicrWS0cU1df+zFTZjHlZ3UYQqCJo5JxYMbgaWWf+Xqeemo
5fNfephNlVbUvFAb4GTN0tbXCBzryuoCjaqXhvMd/lFxWXOD7fp5Sl9RoyNJlZ6WNQyd0Y/Wz+1g
pNrtFvCW0gFHG4JBUzLRLxGS3OdqibiMg6MvSBZOrwB5e2rPmFRj55lY6S2SymOj7f36UVIG9iAj
ilTR9vZ1dQk7UbOQyUM8n/TQtI3QHY17OH2JpbgSGsEy4QPFe4qlo8HTFXu9TwRyUiFdEb1UjcFd
iO3AoyIoUp0M3LyK9BYKhZ6ZvD/69fNb7bSwo349rfGB7I+BApu+L+TAmM5flPnyd1982J9JZZs4
8yWoxCj5xP6BmtXetv7wMkN67m5kv7tt2Suyy8xpidwHSqMfT8qx7GNST2Svs3awcdcqpIR1oVsW
NXw0+fyfuuj0FfmZr4msWsyeDhrGQt3bcvkT2xRdW+m2nXwlasZUOTpvAqVm7R0I+8sHPlksUgPT
Hcrz0aQO6UAmB2ujG86Hkw1/RrC1BZHMaNQPW/W2jZPydR5iKr7OKAs1akVfMD423UevKf/FjjDt
PjKl3c9h2yfRhYP/1HePqPo91AAzwbGxGYWHVgf5RCByBi+igC3E+BnxjUevMptMd7wCOkbKblgU
qXN5u7ESpx2pzuUjnbqaMhT+N5mqIuGduRKCvee+F4Eq+8n3L0xHNrt/ZvoTQi4WFWxtH2+hMHKE
eQyneYj6+zKKDrLWEmv2YQUtJ6UTldP/fuE9/6U6vqY+nNj+ylAY7o/1Y5GjjZpu+rP7XAuT/rM+
2teNw4QeU1lxvw1bgX0EyAt0gwAPil2l8BuPZwPH/+vaD6cOmFN1jSldaqHrC+7QK6ilKkJh7gNG
b55W6UwYoqUPQhmA5SmW+swNcJWuMTeZm0dOEmnkzOfEpXNdB1FEogU6FhqEsCK6YpG8ezduof2D
OVmyThn7fIHGWuFdaCHgM1JivnS+6lvRPTgJVnQJzfT5kaUuyHRZdyMc8WC/hzjxyVSTRq/J+ZGw
wDrYLsbtR5PNshxZ5SL7wFUt1nfTzhFXw7MJGoJIWCuh8XzVeddh8bZ5j/XQ9n7vzkigmPA1pH1K
PhFucmILWqRfKc3kJxl9AUSTZRrRO/SYbmDq4QUX6lyZFdT5vYuWqawZHM9vHnp1dy9CnGqHM6p6
fwKcgRKbXZKiDW03mIAtmOkHLB2DBDF5PqQS73h1GJ3bZ+oWjpofHZMSa04Hwr/FctAjWgJ6Lf9A
qc7mp+po9W4lnQLVMWKuUe9FiqIxxcan6Lkj+JwaDavNJpTU6JXMnL0Pj/PW8ppxq4CNTpOtiWUv
51HL6+WL32JLch0uP49nHKGXTgbt06Ksp2Nc7t3QlXW2QTnoknzvL1Ekjt5rWDJLuEE75Iv5opQU
GEvo4Z3F61bRt6ZudT288k9Ti9e4JXotFSrEXYqqoUG9h24BHsAR3jsp3hSTDqhmemVpPFB5k98K
3MFeKsYfEE3KOS0QkVpuLUzclLe5GWZClIHVDVuJAWOrvXxp/Q8e+x69iO/8B4hGq2DlCP5ygbPI
UHXmlkpKUzBCUn7EVC+2rtyJidUkgSHK88sBupKONpC07ePjR3XQSWkcK2ZOe2Ws1+DBrHLzmPfh
05lAUReAQLlyyEntdPQDV0YhMs4ibPQYBIbaVoxfWeKd7FN/vkwYIWxRzZjplMA1WdHnn56o0TV9
QCqeVU4ae/3INi7iRTgNpqdChd20LcOUEguHa6J3i3KPBzIHU/nAOyeJFjmu6WgomZmbtGQk5bT4
8b5xJEUEA9iXG8ASYp6pd+kofhlG5JLufrarUrbfFWdGweA+j01aH7zHDY0wG3IiIw2isZ5+Scok
LTrEuEvgBIAvlzmwojbT8oefAVepVTUAp7r4JwPP4B9GRXWmld5UTExjqfK+2o/5dvGzMgUtqILn
rKcHtfkqGMKOsNKUe9QtnAiJpsBTL3PsVIcb8NlxmKhZMQF4z3KAeKxuqCuo8DXyu+5mh8rWxpP1
57ll9vix3rNQfgFq4XzlHb6gUpKQxHK0Q/sMNlFhrGc4RGY2wZvxS7raKig8lynYInIf88AYEQHO
EHH+FuoXYY+WwS5TeTv/hX+1AU3+Eun29XXClRUxSFa8kDbs6J6Qh6+K7VGcuN7okVB9Pr0Pxvy1
DifaGqcdZBR+IMA/7t78HiiCiOYfFqqjUWMDO+6n6+4ERnB+mjnnR6/CUcb2dJi4jn49ctXyQkPW
jXTHn7Vj7ADpdS9fJ1TCzvI/LsvyF7SFOSTV6Dj20C/XadVTK7nSMlecdX41nickF1D1utpMLkMu
u4oOKDuwTQOHQSC8KYXBwCETPUbpL/FETU/nJPdCIYe7jA7Qbom58Qfc7piNGsXQ4R8bDNUUMHu3
CH6AuOJRX3iBKRTg3znGytS8qxzsFlutNUOI3sZIoA82rUPYjGv3uRuSvZm9lugVg7WUesszbfp7
QMKQIDnak8KCiEx/Sj/Pp9UpI7qUnGKmTgwb0TRAKjneaRnm9WHUUhktOq17UxWau4lhqJrUb81F
P+Crb+Ht1i+1WJzh4smhXSG3vA/RiBC9QaCAwsfc5kGcP7twidjq2lUtgXACbZaZhYfwutX//Nif
C+2nIGi/IXPgJjXTAjDbVPliNKDvunRNhjVWNRZu6oghjhRy4zSFNooPCekicroy925rzEk/LHC6
HZ4EdpejPqQr2EnmWGoVpfQn5snPMjdkqDgpRiIH6Bjfp6p9opo3OQWf2ly4rne8/r/SmabK3cyY
im53LdEZSl5LRLqplIuNIba+jfbGaHI+3NWf13LlV2RM5HR0JzauETz5SXUNYQrDJgLwvow/yOWg
A/Lp2Y+9WluZkz1lowLGMk6mrX7S/pYx7Dfi0YjKjPSYyn7RKa/U5TnnHteL/F+iwKd3yA4pMPUW
nRiX2Vn0kzLvdldsxKigBjVrvFjtqvDrPX582Rn/I5XKjzmxuS2+1sUPfrVjrAOd/54nqteL6GgT
14NpGwYwcdEyNrbA6ukCD8bHgKn95WkOSPQeV2a0Pogrz8/BNrusM0K5uqenmv9j+n4NeSIeW70I
lTle9o1VyzMdIHEs8U3STNSbn1nljocCFzCzSALY3dlY4tQLk7VVAuBXYhM/285SjpSBursswxb2
aeOTurDzyDhNBZYgLnSSS0ED+RdchnXz5VX6lTceO0Skn124o8QW3VVn7vuj1WBRB2AVNnlRd8FR
lbxKZfFkpsC3d0hrf57xzNLSFG3vpNXs2V3XUaUvN7ermxvLaGPZpXp/xCGfOafLh3VYCt91L0IF
0xYoYk1RoPoLYIyuWtGI7m/w4FE8eAAaqS9s9gQ0WeGCCnzxlt/U74qnOUEazH6dcGB77//w7+/9
SY1vaSSnAqXUlp5nQ/VKlj8yIlJDhtCLsXa1rc6btkoWLF7lxSc8wFWaPh6csaUCPlLysvtlEnYM
UzV24/85Gp+3OxeLAanCpc6dgKENC41RcAwn1Sf71C7FAcOseov/EMhka+7hZMlfSKPADuGZGqZq
SURfr+E1JAfcMbysEieKUlyvJcvhpuRyl5qHWgCufDVi6gnvyVk2jW7DMbk6z0xJZ9hBVamcnMCN
ULn/6+ERPzjwDTae4encej4mRsFNng1Ck64IHsLIcn/GAD4SvPdcX/iSsZobnxssWlQ5QDbmQsom
c0Dybq3zUA66L6bSAZoEgjtnNydiR8soqk9HVRW//BusQGQQlgM6dBK3y2GyyZoGRJoJR8UCYStw
iuqX+NfRiWO2Npx5x+iIU7ODDs2VdkNf9Lp7DILTt42wQHYsJnNWjmPpKEAanF0/iKQh4YdEXk0k
x4cwxlOqnbPH7cJPImrv9tdYezpBVHxyN3+mPXzrUtK7FQ3BSpYiHgHtXdHfiVIw0G1XaN2+aqTG
rtCRrTx5EsSL8nZ+LP07GIQTQtZVLxuLZVW+sWP9lPP0/ZEMyxEyJkT3DhRCSa7AKSk9qw/mByN6
MkkDuuhHd1tiVhqVR+zEaEwqMQ9WzXgyu4SKUB9HDTOYRbuschWjtyT7GcG5l+/uzFC/xAvWWK41
qhkKoG4YVGKa1TIVJICdwvpZbUKRo3oV0oFtJkzZFF6B/4G1ptLPASTtbeuSHTmiSIF6Up03wUN6
ZV6k+NyG3Djf9ZNIQ9tRwNFGe0ohkV/LVgFN6laKgHQj1SnSYw4qd/SddlSQLz4lHXTLz7sBhczI
3/EVBaLNt91UtOtMwj76ZEc3T27sv82JMEpDhUF7OziKwtCt8KL2culrdwWRo0AgKaE2wxL7/a7d
AuA6FxT3IjvMD+dKLOpNS94asK2bxWPHLo5XaSDfM4IFqjSrfdpKQxPlQlmQqYa2af60JdZJEv48
8fpaPDIhyFAJlhEXZE+GuIgNOgctQLGuzEke5p3gZvRj0yMAEn6bwy25zLvKLgaI0mSBkYZOw7nF
5t5xoVQ+qDqDzPsqntP9T4ZAIj8MJZlbhPp3QHQ+8TiThsSoK+kdTaUoef2HYzAf6eX+b9Z35K1m
e/d9UiY+2NEA0GuL1b2fRDt2oabwLMy1qT6JrYb24ko51ap6IlgVB+yb2CA5lDF+1OHbw9z3hXr0
OZEyKfaunEYiq3We4q3Ta8rrUZUhDlg4SH484WOAB8/j2SmPywO0LZDiI0rqlWIDsrvXdBrmZ3Qv
46zWrh5i0ZqkEqJ51gCJdMby0IEAS7zyNdBJNEFIaCgFj0jA7HXh4yDCQimZS7et/wqgnr3QEcW8
sSQ+CVcos/Y/9AoZFzQxhpCKqbW3mpbcMgMpS+kyLJhnU/WT0YU0P/oYZswsipa7TD1QojWNrXeX
af/6p0FoxtNtdfHwoZwM1jire+/xkKiyFMrdedGEQZx94tWHTpjpDiQsZb6OXpjezYau+3dJ1/Dl
6ZPD6F4/Y0mOKZSTAFArAVO5lxRpLr+zQD6v7Kyv6/72jOQe3Um1AZK7nfALHXXG2jScgkVN8s6q
DvW3+itF3gQjWzUeohN6iu4JUDD2pRhcheh/Wypr1VycyQ/VWLBH0aqEUTxmJDltlpN2A8ND7PnN
R3KXSEg4PDA3iKrWsplJxxGx2vfiamTo5+DOcPagmrckze+hmh9wct1punXYpuMb0VmUsp2XE1gD
1Jr2D4Og1qXtcdFqF3qivu6MdjoN2DURKfmx6XlvlAdeW/YhHE00sDjRBnjPGSi1+30A0t/iTT+S
jVRSalfOLC2Rf5agmebiopheWBnl7jX5+2SfE2dmhqzYGoQ/eUS83aTTIQ5qBannugqtu0kcv6sh
9rmrINAAQng3g5yvVrFERxmRcbiWyeMCG6qupkVTP2M6oHiSXWCtZuY7RusYRDGAA2vAK6paFB1b
w7WFM1qEPv5VeiTvgxUhDMnVAO5zUBp+OicxcQGbZx2AWh73qJ3O1LlKhBNpvZau/n3c1NBjkaKA
kL+Fya6o177vVTbUtGiqn0oZk1xyyjFMU+V3OHZCrVbHNVqkkokwhJ7qGwnxWvqo8wYEIOsJXN33
2cHAt/GMD/L4zwY9s5Ic9L+S+hQ1WJwdf8sC6lV0yJoR5P5FeuTUjC6rLhC2bFTT7EPCtBqNOsUP
pBBLR5cpQdc1OLhRgTbkmsrzlemJex+cvIV80czPsDwAiyVEbA9SrWB1u4pn5yM+PEG4SmmMNloB
cPWtuDk2Zq77P03VOUjGx6EIgUy5VuBSkTkIe5WSl83TgEbB6rELmGK28ySki8YdnJ7R7nQGhx4I
IOB0IIUZRrCckZcH7AkyGbV+gNxIzeB/0zVaNN8lIA3u1nDopui7e8pdpuka4c9wDehMEVCCEY7n
L009n9gqLowbtWiwIP97E+Lu+38qv5gafUhG+HBRSM/uv9IT4hcSCDwOn2RfwKOMvJ4z9femkXnb
qDUhvHIV9Su1fULhg6COnOJY02yaPCNZiEBR0JxQ+huDGgfMZjgNPjkkpBGW5noHACJxosv8rbEn
MIz9J3ZPabRHjqxd4VX6ymlyW46RWw6Vn4C7nrP9zU7ilkxLLaGAhEixEeN7+rLncqQXiPbAhQee
htIIYnYTIN2nYXU38GMg2aD5odRnF98LwBGo/C+1Cerb5PBgrhm24RJCO6twXFspCnFFt2fe4r27
Mod4G5o71heA9qIaeRxPoiRJpQANFKALumDOl0wduNZe0QTCwPV1+JIiKaHELLYOxn+js/LZKDCt
i94Bw9qPoT4ObAGU+jJciY1ceaiDNf57M0ehqZDYQpKhzsqPUTgS59Q6dLTQ+/sh5qDAnNjvxLW2
RhgDVQYUWSFOXjqT0XB0CjvvREEhUDoX+m8O4sKe29WKUHJeKZnuvcAJv6p3Mu12ZcUeGf2MCvrV
nEoyZtD1W5ocSnsBpuohJ7TX8kcJr/MBGssOmJXQSMn5ERgELGg1cvvCWIRhjS2P0Xqa0UJoWBO0
mwqVVvCZtgHqoYn74QA4NbObu45kmbWuJ/elNYkUfnKnws2gE/zu1+PQUlYN2U5RkEruDe3+IUsV
cxk7WfqRvN+2hZr3SVRwKH4+ln4HeaGPmhJ3T0GCk+0n6Yeq+GAM45X4AQwXCb+YzEW+3TDEOhCn
ZsCpRFDgOCSKe/hu+7/i2VZQ3p73jWLwcFQWXplXzerijFO6J3/zeFF0RgxCsdhKpkov05+Ak9Fx
d8LaC7kd6M23zOqeQ2xZ+83vmMR8PAgGxcxy9+eZSosby1KzBL1xx8iGVVihN0JZdxobWoOrzrRh
59iKpI6Qg49sDnV+Us6kD9cQgvcXirW3rV518x+y3arOJgmBleH2/l6L2IxcvYSLY6a5kUjLDx9W
7vRr/KKStLVzkbs20LXOQLoLjfvQsE0TosPeAeGNRwjtIf7VX8h/DPrboGuFNPtN5I6ty0w1U5wO
CTlhWT9KSeHt9SQx+g4O46ZzroBscpSHm4tHanVd9oyVQDgkuED9Em9r+K+ECsd1p09VK9n6viYE
2Sm0TZi5uGBZTRJwFCyFF9Uh0O0uI/aIQNvwpRYj+oqLmjHAZpvJsLen1OVjNxbWq/3M4+GSk5P9
pyiZyjH6wcCaXCyZVTPTtCpst+OJRwwQ+QH+Oi3HgjFVnpKdpJPyBXCSnETFR3v0IOkFNUTbAtTW
z06xwNfOmQ6dbQ+Ac7y3VWq+dcCTjWz3W6LOZstPmKyci6EnOC2Jh+xBbnZRqqijegDugulU5ujH
zzeD6HbfVJvuU3s5J2MF8QIRVBasNDs8DlhyICrF88gaMpcVE+c5M3BoWfEVGmi82NofQeb9+pzn
v7ZthGyky/6Tu27+6dYtcIqBt9uRL84p1JMXKxaUF1yQur0/6UYpnYKBtBGaNKIbAufl5t1VQkNz
wM3o++VQ8XVO+ksJuaLeItbYRikrrru8GyGYsGyLwlSiJRIaO+nkypcjacBJ5LMdQHfdQgAaFwLs
aWBHcBf8KjPUzIb0+951DIcizfsBzKoX3UDrZAQUSplY7aI+PbBdujXb2CsKitVeJ695QL00FmTA
0f1RpDboYKPbxbVvBfvM/YTrjRdl9o3cYm7GsmA4RC3rKEQZlNgunVfDk5oM9P1y072elQQA/LuZ
S54g8fORo3pk9hj8a44ub6EX+j3reIWvNZmR6aiQvpK7NEDjPBtRQNO4ppJPOaERa4vDSK+vqwFk
2vEEJ6VCIddUS11TaFBiFes7cSioZNhrknR+EXX9vSumDwN9aQVxvPz+52WonTvxFF7yH1u/IFBh
IzpJyTDkySrVc+VJ8kOF2hjaGBKJf+PHXmHVQGptV0aF5sVChRl4Oh4Y0yBt9NFkoIQoqUldlHjP
H+LLAMVmeVDHHi8Dsg06HLu3tblXMe5j+qeAd5GlTeOwL8hMVVyOsZAlzu6g+jX4ZlVhdwimH3kX
hFN+wzGt0MJSeeUxBs7u5Xn/87saZvouZYeqkc9evUeexIUsojnQP5/w88l7tvYkmvry23xgUnSb
7bqP2BXWOS/OjFaiqXjEeh5f+PsMuJJxW0ZhLJKaMef5gqPEU7Kr9TYtgxu8En2mPt1PZKCpkwZL
rRkqnvJ26GrwEWdzxU/mY59Tw4pBmrcPwX05dtKYq4s8LRIpkm+flbDu+RMhLXUKLz1wf9emCUL1
rBktpd68RYpvXz0PPR4utTKkN/qXRCFONqeATqRP06GJWwIjEeFSXTYID+galRYPiRg8r8idOAkQ
w8wz2Guok2VGKTywNzoxTiqScxpnzAb5BEGPrZdkAAcLgRWy7kM82bBsf6IugIQ3EyM4Xsko4JZy
CU38LNnsEN8uITjxd1WoTYe9xMXbEbW6nfrdS3o2aOUYnMMLyWy8kV1Uo5xT4jcPrDq3595ap1e/
T/kUsDFss8KA5ctjlDAiig63Awkr3gB2gTSHTpm48MWOQpQ5RCNTO8R0fiwdZdm2mEDVTCzT9O5c
BqRItPO+UVXmo+e2pSP/A/tMQCEbOutgfYoJkETx6UG1Pr1sP97qaqajg2kbaQ5Y4NbQDDdAFXAF
D5cpM8uMNyARHI6CMoO501fW807M4tm5bU3iggatzZVJLQkIVvg1mOu2k+qL58TnYacYOdxlspRY
/C/pNMeNWVMzvMIK6DIU+aHMVAEx3W9e6nekDObdjcucYsceyZOkjFl15Aj5jf9zvF1RVYvc8a9x
OaVWdJ6gZ/GqwUAPNebH9QAue3LQLzA1c6ukEp4coDuaYF9zABse5R/0rDYdGgkmCQP4w0oi96c9
PZXCQyRntRloTRszojBMovkD+6KzKXem87NJPvtC2X218xPHwMFO/SbKyqhqSCFWKaE02vJvKBhV
4EYAdFwsOpqWM2uQtfIOkZTGwoA0cd0YWryfQUDQuxBGnCpjfCuSTmKimZgyeQSbRkUQisyOo24x
t/M44vthFm5GP9oFfM1bd67PaY31AhW0pC8wN5ykWooF+Q3Emd/NWjAkrsy7Gv135slOHf1Z3eW/
EfwubvnKWizw8h9SHxvog+Mdujwis8QK36friQPfDTorhZrrQ0FuuBnSm6UBOYGtFsrjsLIBkWcv
KFYIJukMCZ837Mbu0rr4y+2v11eWREQvnAjx5O/ntHd+dyVmwODSioagsTZiTDdq7wJs/QMCd9jI
cFViJUgjQ2XYbeiCmACePAR0IP3dVBJDXHCmyc/Ni8FSTttQ6DfOnbQ+Vzw/p4H66uFfddbw65uk
MxZaxGQhRxkPqGoLciwGNHDJYXlklWiE2z5Cze/snc8fae4GpJlgVuy1V1Uu445gk1bXM6CW9r3e
9DznNnPTsgWbJZ5g7Mj9w0hpHt6TPuzrkAgSCFlksdVUTBw8pXR7cATZvEl0iGT+FoqThufglcnl
3jWi+EE6AgpwNDOmq5OR0EeH+RoFpywGOhdUOnityziaNK+opSBt5LZ/VOEGFL+SbB9xgAGZDpJC
+DqHBVzXmAQFNRsM22Xlzjhh4Yu1PwKO4r/2CH+rItf8JfroRagu4unTeUz02dSz8o3ElRWWUepw
kNHX74Emoq9gKvpLVC9t+Re0wTTyjENZybzBr7UjdPuXK44PloJCeog0yJj+dJ8HxVjzF0nQtFEy
Xwzy0dxhvE6USjlu4WRk5k40qowCWcbtStdobAREJF+asSwSeVEmhDh7lm++nIfthVCtVqD/Qo0m
Semzujish8wvODY0a2PWECsJ8ysq8UUcWpcesR1kPfITlRZ6/1X+Ddevq778Bj03gFAh25y7zVN+
2uEoeG1oNdynos0YPpdpqpYUV7v3mE20OED67+x0bjhrGQFx73vdY1rsXV8KnTXaOnSuSQzmD5hd
JPghMVcrA4qUhSmk+Xr08ZxnsNxPOETgvmJ/9lvpRpkipMmjCzlFTwhOLoBYAc+R1JGNuaBoByID
XJ4523b8UGZEueUmEEbDmbA7xlzqphh85Tw4AMKwI8suPSpTSyvwPpr+d+AAiCTLYwTqmtvo1t0y
4jJvf8VP/QxF/IoAj8Wp5hQ/WcMwKwMZq2jj5UfSGWcbbPMvZM7FMwmSpYLEdAqLYeW+LRk9XmgJ
1H29ALzkN5La8orDZBd3V4oL99SSrKcPVwGw0XWH8UuKfN/sGApOvkL/MPMCe1aKQ8tlRtIm9UG6
cBAGt5jhR4MA3Qegu7lR6DYE7WN6OCnl/nTOf83096BhuOaqUvhBcn7IUvsXDYbckvkfNCDFzCnU
1At88DLMw7q8AVfqoWm/SuJDAMPTVKIfvyWPWxHwiqi7XFKCLDv3+g3bQDRmoKGm2h/bxvcQ3Qd0
DGOpw9MeD3klfz/2+1m8VuK4YtBX+OtJcug4CXSebErJvOiiLkCmf7lUq3kTCmk9o7b9rlL/4DLE
xIq5fsFkZaTL/I2660DDvS5q5mat52gALKPDakLcBhnUII4y1xqvRbNB59vrLa9N1nzosorsJ008
Tz8F02mwBoUoBfqZ/8l6A78QmlyoO7MDqcyFe7iJ5lUr9Fy4BwnFC0J1DkZBdqfbVviTy9r18lDJ
KZ9ip000K+56Ni2+r9AoMzp5RFdbaIoxyMnRy3b0EJFtSMAKm+xrvntupjZCkAEh1qvtxsUBlaEP
otdzyQ0trg7WD+Ugjr8oypYlvIshaE+vNPFoFq+BjM/UK1gZg/yJEQt0bPd7u9WuIH+oBzVx9N28
V8pO4Y2EnkR56XAse+y+Fk6eg2+FeWcPmYdcF49RkKNzLudvMw68No7d6ylsLdyW6TdrNv1AR9z9
eP9c+Ll3i0Fk3m07iszS8wVdkx4JjwuwmibTTSIMdoHW8T92Sj8FXB+RgddqAXMDBxDlJPgF98Bx
chBhRV86kjDKfxmY5lsrT0Zxg4WOHwbo48i+MP44M1dui6iAKyLYW6ouCZ8bNqRnWefNPnW/OLIa
zhIFXv0nmG/SscFCtBrksW+BBoxzzVQwLZasGG/St9Y3LJCDf112yGubR9I6ZaqKWtJGN4mYpDID
0QvecajP0KGq5PaWOAyhQsKwWESBR4Im43nouI5j3aEP6tF7P+TsaPvrPrdod5eqLzylJxgmdVbr
dA8TE/Vk3w4pL5z4eyRF9fisvtyZX2VUwP8K5KBduwJsyx8zrz/2RTZMDUj1k6D//4++5rLpRf5h
zh2lCLpQdn7gM4qEsYLsy3nH7AASxrh9fbjmmFdVD77ZLgTRZeBcRpcWD1fnqQdriQOd8Oi3WDvu
Y2EutH8pt48ANMWPu+rTO4Gu0u4WfTsQRPwekoaHlDhQzQSKZxg5Bbp1zy/fFvoSIyhb3rWW6vQ/
T0aa5lYSSoUK36MVC7Er5gINpm4So3L3QkaLo2A56BXj53qDhCUA12T3Twe38ohJH+eijoUd1X6V
wnNfAibWsJp9+bS+2v31FckNHiZvTnnuAC6yvyvknWo6yCpkyoQZYNQkOCMPcJDLKPOKB6uT6N1a
HahIChFKFTL/olb6A3AAVsvXhHoG7OTd3UBwApSyqlY7q9NJC+k9WR9tPMUDRtnP8bo1jwHRRexe
zNwIeBIjMzFb21DSkDjjP6lN42K1mwTqbTksrPLoR4+D1Hby4nKclCmFFDZDQC92Pa6TPrtH9TII
Py/0Fp6vepQiXDVHAExJO5aRbBySPZFy4f+h11r3gMid6YNxf9jRIJWoDCiSTTYBsK+9xrdfHZKu
1Wwq7Lla2pHmiWNxQ5OZqoLhZu4pRLVGF4YuFiDJhbPfDrHFtnetg0o9vyM3Bs2q7V8flS9PaQXT
X0QSeX/rWCr4SwfDDJ4e23JPYGH4PVoq4sK3WsXcpFJ0MSVgWnsTZ9sMdHoIM6DkLhfEBj+LCadB
aP3SqUIGeQ3MuJdIuWxzbpcnWyawshbPlAxROEw+H7L7OFLy3FYlghMikT1DLMLKkzq30BCnKuB9
7ijNFa1ltC/H/0rcDhUf5is7b4PofkYh1pCPuPmGioj1P+NznsnWTV6uCMDAaBt/ktRIRhZXfwJi
CJQy+Hy5AcJuHJMPDdgkvYk/W2ViLJZ47nkMxQPvaWdHQFoBMX8Mj+YKC3sNpHotmdNiWiYkKqHy
KJjv3SwBXBErbaIG+4elI3yP2+Dhs9p/Z4dIUQnzNRNkzOQ5jBkVAUpegl53kdeUpv8Yu1VHhgeZ
/IEFGB67MGYcR7pO/r/QQMDBj6w4DLArv0M3IUhwmjYDrCa73Eo7XSJ0e5UMP55do+22qHgHcsYz
cOBk/KvFrHZ/lqsElyONRRlaa/hlT/ChjguSr4Wepk6PlB40fNWhJ62BKtzeN9mUquqXikvxg+SP
kmnvB+FCJkUh+SRqrmfbk74QVidEOVXRAqRXFdQv+JrNdRJHOYo8Vk3CESkWaLsZjyVufF2i/Nbj
psR0Qd3MTklbVXAYGILrFRb5tdvVCYmE9dVss1UhK9wrd2C4P61Wz7yH8U/cWQ7DnOEZFFbXYFO8
WQ0R4vODhZLCbf5sD2BcgXAogu6H3AWIhdeK4yXrnz2vst6PdF/YuBoX78R9ooOPfXgfNJ1GTn2a
40iW9GvvQQ98n9ss2BA8DF7w3HPU8BmgmsJ6fWt6P+w0u1sQ4BWIv17CcB9hT67lD+dcTlXZVfGf
r/GwueP7e4ueq3ojKu+HAW36Gu9XUJ41Z0XO0X8OJXXUeV40iiONE5uZJRgyAJRMrJ4mWZFdeV9p
l4aYNB5P1I1AkmiV9bVPYeNv2Inn2rM9hNWpUf/H3L1g/ndO0+aAWtPH8MAalaKg1L4CUTYNNrd9
EOFz0GQ2o7YT7FN/5TwJrvjouf5P10vY8ExBi0FhEkOX8UOeCb38ZdbhcqqRTVBG/WXUyeDhpaGl
IrEXSZ3WE2QLtjIaJPeKk0NfMMrSJzzD00GMgHh87WaB4Zr/GO1VF4SGKnOHAOua1HAd5xc2ewqo
8k1lOy3r6WXxaAQqcgG0h3JoJMzqRsYaJi+b4cNpMJGS9ppS1HEudScmj0Vq9KM9MWLdLoAkb/kO
iHkM5YaO/agmHSGrGJpq5+rC1WeADROn9iowpiMOxmuZSpcC14RqTRJO8oD61gJ1+iwcjtjowW5m
GWLTOJbDeeOkqQ+catApsf3kayBQfQTIB1kfiO8wSxR6qGqUq24+dsCTmeK/2H1naY9G4JHLzuxN
5219HD0GVLAJc6SymXki9XiFMr+KEn2Et0IIJ5lc0cZ9edsV0hlkfHgm8rTLxtijWCoKMlqC2/3X
qRxWZRGsZ7ejBo6p93TjCeWRfi07kejGfA95cdeXvjNrMBXJ3qMER2peCJGeoyDrJkufmmoBeBFX
yZOCxFFYih9zNhCcSaP7C2IX4TQja90pxbLeW7V+pNtVbDkIk4ZkcJTCFB7MGZuMEWDsI5vecK0U
NN/LlPOQPvkRpTWeePQ+2KeDeWr2AHUhlelxJoyUPak42Rh3gcgVFQDjEdWJej4MpzvHmbQU/Aw2
rKw3AbY6yd7lulB7TsbYcbqrRG9deJ4WM40V9XKJcfegOwAFI5mrBSxnhZDjw86PwHrR2/VkyeC8
ejH/Tk/IUdw/m1J1A4NtLnnt6aZtXLwY+aNEq7i6CSn9MkklRWzDIa/rksgC5Xoh1XeHZABUSWo1
gDPo2FyPgUOR0+ryGSW01eBtH8E9hoH9PUaJ3EzlwR7x1EYxAy/M5/emUxoB+SacZARTo37GzYck
Ja6qBEjIS/ADI9Qu8JYIVZ5ysn7MI/O10LV/xoWJ6OwN9ynJBwc53iv+/Xc6rZTZkaHw76gYH2Nm
+rpZIjcikCL1Tt/3GU9qRNjyA3H+qOkOspOJrePLRq10GUIHVFbyUiKdUPTabZKxiqM2xW6DFdKt
hlvc9eggaXmyyHncquRJjljNT3mxGARs/lJHoDKvTx7lZqyu9MmVNkFuJRJmOZtBaKH5ih0nnEFo
ALSGcgKbX0omGtRwvpHZv5LIroGS9TdNZa12Rq+GUdVnknMSpRitqqiOOPE+hcIkLffrjmD2LT4J
q532k2RNzUWzGMmiWaYOD5kikJ7oc+1wO/7NGRKdgqAQuGhNdS6Y1syhUtkuND8/61X8OcpNeclJ
vhE/H/T4XQPU61AS82ryBOOiO9kVw8Td5HEgBHn7AdoEnmDnOlWopBa31LBPw41v/B2Np1xP8AyG
ID014r9BImPaRo/QgvJ5Jnk6naWviuhsdlesLL4S4L9K6DRNu5Ya207783vzJ7RwEej0rUU0dwgZ
LfAyRkAdQOhp8kjFfZRckQYq9vc4IPgm/IKvysnyqZ4dbEauu02JWWIBZS9SGlyuHHc3jVPvnU7G
dlG2mFSdaXTEoQaPWb2Mw6Bau+aE8HFPyyYan8C2X6w9likTrxfAd/vBi05pJ24BMx9HLcY4Pt8r
ShE1PgCBHI2FvZhm2z2/VkGyVLbWTI8fadriK+W6K+m4DRIX4Y7cyeJQz2chKa4H8vyqeDuW6YnS
TKmFMX5+G2pVoZUrOsLnXPRmZv9ubLnjLWqqIApLHoMO9eOHUopK2lroiUiOVFisyTD87SWfi+Cj
hIKgqCsCRBr218wDben3JYMhy3jAT25V6Crj0akoQ1SY0uvLNAc0V39oO5W2YkVqfnACXQaJ5DJS
TDe0jpCunuwt9BSKQ2q07tkg3mhrvzgYIvukDKDr9DkyzLfEB+hJbNWwOrajSDXW7tffN4uZ+KCx
d6hOcWYxiCaJj2ZVPgH8eaXgAE2mJjlyMrC871iO9SB0mJYKIwRajhRBwl9zowbqF6P5NSHfrxkI
u5IJ1RIAnTxK6ye79ba0E9rxPDQCmSTMFWWMn/n3Ix3GMbeJYoOFyC1+am/+GQhVZkXc26HDVtxk
ee2P3BnO0miaysEO34Xt9Mk6LONFN4JtP4n+Fhdy7ko6vjUxdF0i1hsprnirrFeoEr9qP+eoG3OM
m3CvLr/WGo1NkzbKAp+qxzqQ+P4DN5JMYhv0wLDyDdzXeHdJ0syX9I6bBQcAE0T4RuzZmYfrW7I+
eiAdvu5chTenteeFa95b3s/p1lXb3go/b0GQoEg8wLJja0YELtZLMYFedk8eiS+RdwQ+JNBU51EW
vGMBDD2DTXe0A99jLJuSF9qlgLfIIwRj37bOsrJMC9jMJCO8WWDpPpCFOn+NqBRaUstv4dZRFEXZ
vCaXfrkdetCk1ZHyrrJkUhxCHJcOqDrRoUT1a7EH+Vyey7kSoCU8alPvZ7r3+4V1kHTtSXokFz0i
YMjZiz72yftBTm4on+I32nFH9RBr1EoMU2mI74w7aZVmo50Lck1Q5senHNKIq647A3+r/pnHKiqJ
2suClyqvdlsRojsLDkJa5TL0eOHn98LMG92/LMcUZhKm4Yl5d14lYLjGzrZtyqMgjGIfwBeeZTOS
/4uffR/FwlE5DOn2mdn5nTpWnt56TP4YxuRP9/IRCW5cSN//Qik33rsoawT73SCsTK36Hxa2WAqw
uzUsQXj+SWz/9iRydeaAxHWcTNuuzI62TuWw7WGwHFgMlWIZqUQDgHv3RP67TnV9cKv5OkkkpL3O
dzw0valfFlE6+IaO9KzsTlFxA579dPgbD3Gv2DN6iqyAgBkwjVixqAgn807O5HKseMw5sxOcbnYG
f4d1avF3JsZYkzMQ0Jv+KqFDvfMaEgBo89yM+0Wupk1c2yJc0CjZapvzggFLM/uEjOVO+TD2GJqk
Fu3WfXjwRZTA3NuculXiHhrHT2QUtKBBaCrVEWXT5SEvtkl45A4kNQ71oUlrhSasgzLs7rKIMP8x
0CxQMWwJl6kr/+l7ixEzsoBxzMuHgns0e9M2UCbxcY5T8/NT1391K3X6IWy2hRtirnGrUPrq4VCE
EaRheHICOZbbh6hY41elcELjbLJIi/8EJvMxs7HcPEBO2ahp5Cj3zyIh3d8VhJ8cX1LK/vLt3eSF
GtsNYutzkmCY27LOPP1RFjROu9+UOrP2p52n1rXs5SQ/USiwaLfj28WcteYvlO2RU6E6GCMIbodv
OOg4Jx+9sdcXcXo3eTV4gjHaqYUZVhR+aHnU/zRzfASIR3b6S5xmlyJ3mptM9u6bnqw+Biy9dH/M
HbnNP8Y0w1yX389AGddAV0vF/u0Ych6XprvqPrM9xflg/bEFFyOL8b/VXDeOcElodRpE6kqKTsm1
G2gcxxN7jjhSllNWDgEzsEU/mEoydpJiwWoYTzPeSz68jVwlfN0z3gzu5MIAIhKMB8OgsVbYU8TC
8DsdM8cxbUSUvLHUhSl3304znZtj/v6qj1YBfz3Wv9+Tu33UNjwswsVYaKc+ql3GtJ4zgolsFH6C
SR9okVj3LpEmWNf465ZIcf2XIj94HTzi3XkX9I4hrUx9PbTNGk6Z+ja8k6fHKjkiXVEk94sRxVE5
jJZwZB8hMR8IX4KExVyiUr6MdNnoPqxQI9R7q7e1FFvpaY+kewF2zukYHMSQjERzT3jgyqrCInXU
IeIlunODMHkLNxcE58AUj+QXYawL26n7r0WHqJyIfbAQfSldWa6dj9ouloIMgIBbkSUBbD2ecXhM
kVc+ongN/BjMeVQetWzU1XxxaWByuyIpXyxkJnW7f0XtLU+3+SkE6NVs5IVf4zTSQGTCa/8JDobP
8CA0WTNnQ+nBnoRM+WCqRDsi3Vi5ZG58YgONPV1lpcS9+3bzpf6iLEih2iExYOXkzQN4hZIfXDKr
uuv2wIqaAuvIQM/TuzSqPadgLYwbJ3+mM3ZnJwmMOjZ2JDYvbU7PfJKYZo+DQOnWsWfD5LsUo59z
oEarwk6GLx6GSYGNn7/pfN44ORJNl+rXANVGwZBiEqjC1TT+1xHC3XRtReAGWUTiAZH+FYn5zPdI
TP6clra286L/35Ic3hSoUMKx/rQaJMyj3jD8AqKA79dnnYf2YOY1Hjfwggxu3ZG7sCgQTFbYAds+
COTeFlQx83ik7KahFpzMYw6qBr2W4t8wo6euIVSb5UINDJ7HSduqUwG+o3uTaYybrwarlZgyHDNL
0sUu/Hc0Db/3xuAlN7qQZacxJ2LKcDnPVFmG+wH+yNRxPje//oVn6UE4kxu+w7BMbCD+a4a3Z+8F
g3Z1henNIg388DYJ/8apBKRxRKjql51FRDknNbmjjIV7tdaOtPEowhgh48XTANaMTboglImdgyFz
wsTRqdQ8wTrqKoKr+o1II/m8Kvk8ueVRwiUKjbYBgg3bezEJuhKTt2of8dZbaUSfopHNFRmJ8G/H
qmpxsem3kYTRKgXHDBaByy4x+QYSMXZ3i+4n6c6XMYjcVMQpkAe7hWlj9CjWmMGa8W+N4G0AzePp
li8asrVg2DYq2K6xCfe48GYwSRi3k8bi5Uf7y5VA9nVDmKEwHWVgRyGMeFXnx7mScudCodqfE4Ts
10+bPkFe90NuMbAGQOktlHG4Ic+n6RJT/56jUF0niVUXdf41XFDYj31qhoDSyEskWg45VkFWc58K
DQSyDIE5HvPzGxNeVAgOO/uvZMUurkUUbhJH0/+ULNzj1/4NIkPbSd0L9KT3+LNP5B/WDlIbluzW
VODifb/9/7HunzlQXpgFVlZGJqLAuZer2Rw5zcK9AIxjEpf4L1UxTdn2fMs1hqRoRq59/GJYANg2
cb3SyPgtyCVNXQH7ZxoxyzNPDQ76vFXZsXbseXOrpN+l/in5j/dIvC9W15oBdJC6AWgZ893Zq0uV
9tp+PoXFiFUCDBg35J+fkGeKP+7JNssAX5j48Ae3s+KzXIQZ+UxeOjTGiuOPWRdMDUyHsP53Y9Hs
4ZhsseQABb2/IIju81CTsM7n3Pm0jf0SCHIovvroP7AWYA5YjYSfbzHUEttCdSh/4fEnBMyRqwxD
8Q10917V6wMvdfeJljFPaAyytSuaPG25KevqeDGGVdlUxD49wKmeTRmOOiX7OYRswyegMVY0NXZs
mWJZOisPTp+I/7hy9hQYU9wU3X93UcvwXduDb+Bc3dG06bXvypTXSYCpSoKftecIYPQidVwtG5vt
dQkUqbXNWoJYj6DLKJOUeRz3dVWWiTqWHKQAjfwwB6OBIpEuTXP8wrNzkJW7QXpMOaMk0yjyqLz4
TkAD7XFrHdbCkX8SF9v6NLSeNMazd2nOUpsHen46gQMeIVnTFVl7rG1zf/0oHu/emfxCDu0XudFV
uqhJ1G+966sJtRIX0ynyl2hXi1NXz+TsodbCtbPRpzche3jsZ4hr/UAubHkUNvND09mSeovEwDkU
5y9MKHqBm9D1oCX/wO8fddozYQ8ILSxfjZrT+VVNaLrWkmt38wtB9xzAW0oS47DMblT6AbELWPUh
GEaLdcUFOW/Kxqi6SI2qldYa8cZdYrh8S8ayYHtriF4CeHCV7E2AzMMho1Mt8Pmz2IKC3DmIxhMR
Hgsam+qwGrW89AE3mYBxreKFgiL8AnUl7YzEgn+PMZn81e/xXI1FovrTRoMA5N7N2RKX802fx0Yz
Mb8hA7ZsQYILKeBMJ6fbwr78CVv/xR0ARA9aYx6y9Ep5jdAgXGmMExww/iYW6I4dl/BUsk2Tzi8b
j4cFeGvSl/B7NhtU8vYUpcY4fMvuQB2gH0WFo2tj3yWiMMXLOSjgzcXbGqLzWo6DGGOjZhuGPrrO
clWZVb33+z+XhQ0Q+m/KLWLoPqkgVHn1nw6ai671uFlX++dW+CeSuILpoSr5JO5jLJZUH7F4brN1
QrhZvMfGrQQYoIbGQ0DlUiUDXZtJi9btI25d/+8EJkM9fQC/qOnVDhpxVpUybFXRtenR1CQXsryJ
3RuF7LmYMiLwtbiDZZGAlmm+lAVPuLfytrVvxVAUfPNi5pQT5fGjW61IOraZru8FVlGFnEYSiRov
5mVvGhx/g/OnhLRnJSs/5aRpcCZiWvItp8PaVNOjWSJTmjrRBUtQ16WMvRn6rRbX8YNTLOUvGkqD
7aWNrgIoCBrSulZMGDASVLXhvHETHOK9AjowGlpennPYtx02OFw40ucawmxGiKJ4uS072Sxf4E10
5/6xGwKGVHpwPx+ARakmzquT3Qr1Eq/B56q8QzUE3wghWgVn1Td4Bwofh/ugzcP9RUnSVRcWOVR4
RjXXOmDH4o5pr6dkKZ/56JQQKXzyW6817jkGNS+ZOw1PZ4MKCvbXmmi2uAitN4BpUwqkaqJfwxOB
jhZ7Q0qoJ3Xv7dWawlKB2sLDdICZv0MNsMN7LYfDOW3ebzYzQpG5p7JXl4e2KjzuTQpJDZtwUn4T
PKdZxDfCFerpB2N0bS34gD9VhuvRDvu/rnCBALNRUIECNT2B+Z9BkLZ3WRd99TU9Rpz+ngZ4H9yt
zs+Yp84LRSLFApchbNg3mrfqy8h/8n4b+RAaNG3Ef66UJMX4Fl1WW0HjeYZcU/9LSFic/ZPIW54J
yw5d7F87cFjJ4O8rkrFrXwZei+MK2di0EpXClgaYk5cTjMnhH5HCIBqDMW26DeuXnEGMYf7JQ32Q
zOBnenL0CwgOo8H8JJv7Z4G+0Wq272I61+eZCi8oBQ3MaNR8nj7WmFGa5Rc683LV9PiBlxq2/Ju+
fKaho7VtZDlDfVadfR+NieuFaJfX7fXzsqCzUym+fWvJMJLCKpLUixVPSTBOW5sldpXq6PfPk30C
b4nD5/eBfC6JWTVyuu/lBIhJ5Iofk23jju4DFF6+R5wEkV76EykckWHPM66yzmRux4EQbCnnYTZE
VRaiZ3bNol5FHSPqa7hrPf5nX1cHaaj004PuCDM+y0SOv/u1aTs9WoctGvxyQLhhyyF1Qb2twO6N
k2tX1u4R1ov1ZV4SA0+fuN7WyOPHC3epQ7J2NAnCQrigq4F6NHAoQ3tzrHlqtvPRcbQEN0sVhyzP
Dlxc/I/BQrcDuqybOKAHIurbAM5/x+GxML3bbNSK7WMmX0Xc9Oe/b63p+lLHj77zO0JLmugjQkib
9wxx9O7zWB3aHt53IOuRBpETBDrT2HgaMfR88wWnE1nacs7DQyX4MGwiUpOZWTLMa1mk6z4IqTdM
9rBbfV3lsc+Ga1HPJKfDziiaDtx+f/3OqS3QxwG5XqJTm/a7pnCw8Qss+YmAeFHTVhdijl9dN+GJ
wLk/0InccnuEWML1HuARtNRFKi3cIIVXml31pv8qsdeFqeivOpt36SsY8wHT7fcqKW+LXuxqa6Me
3gpZZ6yaQ5i30nhRR4m6OK1jvIvYZdVdrg+s/U6U36LkXErLAN66ubzSwlopRhmYI4DT5Lokulbi
p04m+CtELFTybxcP3HF1wQ5bBSwheVLd3eZBzKqUl9DRsiB1V7KPLaNZIPd4byfW39VbWZdkkbIm
YSAnC/vwNwjeVyjMG4f6TKK9yFL07dzeXBmFqcJVRGIz2sLp+RBV18AxyiguiElUMfcFMyd9d+/4
T9/C1RDWZUcVSweFfZFlHV2+opdF2R+Ahn6IohwZ+yo8XJFmdZvxvq3ITWEIZwCi7lGojvHKVv/Y
Ws5UoSPqB+QCoLuWgoo0Kw5v1nhAJB4VIBM/g13vCds2EtslbM7OBxUYPzVOVgWzbdoUKG8bM/D3
F/qSMCjjKO/EkiVU0/cscjs26dV6HPfEZy8hXsDg4qyGxRUsUKP8cwcvmY7rj6V8IpQBZK5++xSW
qQj0CGn/LtOJ/vmsOUGGwYPwW1QWdR3LfaI3elZ3c5h8slLQX8P3V1k/9K68uVT73uRCKOvHS48O
bjh7Qf2RAc3eoO88I9rsgwAW0h88lit0m3KsGI/iqizUXuH2rAqb7geopZkS8p1FHQRmqaIPH82Q
I/z4eo0en9gd2ElL7h8Efo0Kszoy2818u8bR/Ri/uFBZY74KlhfrTwy6t2RbE9FT0uszz8kqn0aD
WKVl66jgUsgsu6mMoRKsp+S10rzfhgnBs77sA4UV22bu169FCjq4hedtLtzwsj74yAZUXx2OCw7N
MA4JPy5/UL1GGZ49+J6jQWBEQXJNM1kvsFMqZQYH9Fy7zvll4LOvquEWpu64EkUGzbZrqlbyAQUC
fKH0ZAmybDAE59afDsdMHSPZpzPUNcCChHcYOSThPWqFRp0UkxR7OhRoeZmjceWQHtAGdD0rqtIY
5CojvayRHVyvdMI03LNVhYihKsJhLJTIYRuMn5XywI2Vp4PoUJteMmSykS5V8z2SlLc+y5Te+CED
sLF8PMUq512wwiFB7ZKT/iExZoXghx97J8NwO4h7i/wi1ImHLuWN/sHBvAZZ6ReekGz36aGPRHAX
QDGvWrHTMve+ra25sgyK9ErN4ijtfgp+6PcAVWliJDxSrzzhJaO+N/xRkaAQNDzqbjhrfS5QYVhT
RZgliaggN4iiDP8vRJ/t30S0U62snBVXLQuhM5cEXHPfrGmqovSpu4lQAEsx15BSWddVHGyL6efI
ConRn5/V+JmiSZrrVlbddq4X8epU3HFgIeMhkwP7kDkDTukX14qG+wIeeY2f7b1/qvVLTlt/usqs
IKOf/I1IF47/NdRHcq3WA+S2XCa5y2DgR8kZTZCQOb5Hj9NM02FD54Sv+mWAHNdFjURjyInVee2T
HOzb9oyHATm8+xgCekJM64tovMl7mrJhpggDYFyEsy0u2lcaPFvl2cOIisguCyU4VZElzPVrZuRP
MOUMNFf1m1X6ffEYfgDSoWC544JLH1NEJtIGCzqs14AXpDwPUYercpYTe6oOMeIhbjKedhc60dnT
LRwGe1gCGEKvJT2KQeYj94DKyXvzCV4xUDCaYHX+n2+2Bi7YR+Cx1q3pbF/WWBfJCN5AgVEZSkoE
ioOQV24dd0rB286MVK9wUBfVws6xsF+Xp1Wi1FcZOopbSXjsuRiMCcWHPglxEki9mZ59ijhx5HKv
l7f+YHxV5MLkrXYhuktRaEjA8cM/ZYxhWVgOdxIbftIWHTUC99+W60Nj89EWjMc0s5gqDd8V1wTI
IOWiJXHBKdcb+r22DUOF9vqmorVTue2kf7G7oTurMqttxvLNNUrADWUvApMhMI4hekA0MAbrr5Ls
6BaEXfT01rEeNUKMgUOmRvFKPgo8HguZvh0m533FSUeiYPshjdCwq+2YQJQu7D3AhOH8jGZ7b6yV
hZnOTnhEbT/uH0b4nMKcCNlPEs+iyRoMv5Csm2VhYxZ7G42LkU+iL0GJokYkBG4mesgDLdDMFjbq
ra4fil/kxh+btbDodRiWEYekIMSR7mCZRObtiRccsOBv56edkxPTAaXZNJ4U45v1FIBzZELjj1+g
R6pGE1XAr1dmE8NKqrI+7rRO7g6OkVepE3UFlfxNctggt909F/zN6iZs/YD20xmqd4HUV+icw2e0
7PLhNklDS5q693XZaKv022P+uGmuRdfdB7xxVAfYn0Ne1R1xXT0LrMt+C1wbPJ0NwQ85r3Tf2M6x
pTbzpptUpb3p2qZHf+VHXHvhEZZ/Ia4O7pG1WZTmYB4uTrZdrERY9Hckp9qZmN0InfgdbMt9RJCr
nO9954ULQxrOAieJNK4O6cJQO+HA+uziz0AmtddtEKCXemEOYeDfDzML82/bsZ52zNSbiA/MkYw6
8W9+CCZaQk64ViUgxLCRQKcyNaw9AR/hDdF08i7rp/KUJMUl748xvuM9yuB26pcbkpN60qfF/43G
BOERYuqBwu9RLz0I7OHw3gIsbN/+6cNN3839A4leMajBUPGvuTNx5ZHCdgkrSWw/whojCFcfk6L/
qO5hR+7PzwBCvaxb6zkHbH9NV472xcUwPPFMESK42ri6R5kFdCwzpV5LIaWp7Q0BkW+r/SJdrVGF
8cLoeTWVXjzPaQzMo/SwPj/cLfQmEY27Wu4jEgRPeFvf/lIZKn/MTwsAuzrZqjRdsr5lCmGWkMIy
RDzQ2oc6CQenzTUtChCfVoXN/wPMidAfLaJvMImlIGxNVF6Fw9GLk4lhkoh8FQ/TrqCL6FzqIJ3Z
XZ+L6o73UuBDrTzwsp0AKgxMN3nRJC9QhuS0Pow4RSGCyzrAoDMnuX0IuWCMoBr+ihgdikhNtvUn
K9kKB3u7YY4Yg+6EGKZcBlGuqnE6BzGy9MHVMZ2YeVGZ1qRkHUJ2YKDUOkkVG0G4+05DGnXQTKHy
oDg5IyFcK/tmIQiXbnF/s6c1k+ad9mWjHWyP2REZa23DPm7DSVMXf73XiDmFat+nEZIjkBgD7+4G
i0C/BOUavKPJxEs98WyWyOkewj5FHtN1w4BaRR8+JUucuUayxqQ/dLEoHFsJZ4/y46EUo/Q7jp/w
oZ637MPlgVgFhTzSnKTay/zYa1sg2VdQc5vRVeIXxjCfR5lsmIggsJvtM57HEvvsWkuEuiv28kgI
cONT8mhukJtbHTinMKr/kyHJeN6RETvNIiLPoSi+J+CMPi7ImCu0GeGH8ISgfrp5zl/ZUMsQU1lL
hwDJzrGUNYub26SgdM8uoV/ybp2OnUusIjRBhPNKhj171Ez5dDwJstKlpA4XxkRrKNlNk97+LuYp
+gub4vD7kDjPpJXCpyouBeQfZ41NJ5KH2VTnHQRVq04F7BXfEJZFp0Zc84Dil/JOH8YrVw7dORjR
jFeLXg1kDJk+D0YNvfWBOW4y0e80NDd35M45WebGDVmUsK3zD/psMZFyVTBa5eEc+O9YhRaG1sbE
WOzHQu98AvjGdD/ZwmOUq6ULed6iaKqy/813wg/Dkk2YsrQ6X4zYIkvydG7XlOAe8BBjnFAEaW2m
4PZvcP+z76qC4h5v0pedux6O94lBgo5/fOOtJCNUlLnGIxSvwb3oB8B5+tmRRZ0hwVMP9r3s/7g2
xbW42NxhB9mCStv6Rg7/4q4GXJgdOr2Od3EvOacFubAxK2jx0VBUzfAwDc3hl9DX1gkSJH0KC+l9
pOWIcVJ/Li0Pk0gFzTPz0LbMMHE5ZNgwVscj/c9N9kTgLRWyQ/AU3nN4Sa37/bt5inFXQdm8y/vD
1H5zbRI2NG26nhq8VXoMRyrEEXSbiBmmdU3r050sNUEjHek0VRzj8o4rKm0AGUipjU8vDkHBXo6k
HBBeKlyA+vq52oDXNbTaPO+pHExrFck3q52lwM0sAWxUKTTbnJdh9Dq6IZodD1v4u6B3DKNLFqDI
w1p4iek7onXYYvil+yjxKlOGliWhlwGaFVQPryPxK/e5lcMl+92f3LYPDhbfZrDKtYiXXKamwD5M
JFfDMQ8Kdd8ZZMdTW9oka0HsaLtDyAxz1xcpw7kece8jtclNczP8RbMVSicX1SbDz028UGdUzF/N
18kP9XDI/zFjC35HO+PKSIiaNRDbOiXNcVcnFyM+veREZXyjb7OWIX1bEjIRQZd4qfSnFIY8RXMl
cvVU39E/pnO00sNl7I1xvucDzH3+rcNg/dz9RtG8dHEsAZ1JXsgVQ8hwmEMK26RwoDe8GOEuQEIt
jKT5ANcXtGPcHBb9iwaqtPfHDwmodNiStq8Vf1tQ25lz8eCkP1MftOsUnkmxr7CoUw/7iJnJkOnh
EjkrGlj8qHC4WecG/958cUGaDLVmalWYQmZ8c2R41p32zCxSY73wVmLO1XgzRJa/0QMTx1GiLR2q
M6tCKjH5Ff7oM2b3QwTqdbrJ6qMQhGgXFs4XGPQ+CcSkNXTv7C1lUP3kGgMUKtfPntfx0I/rzYjm
+IfRK1HXtqULi+catji68Eo2Xw1FgKA9kjWgIM0nH7X2k4ViiKrSsT5pZOttaRCZRwtB0GL2uIbX
WGWsFmvllCdk3loTxYSb/1ztyYrmphZuuTDmIsJcJHGiMzWS4I+QN5NvK6him+VivovhKqtAfxek
EsQNHiXe5WPKj2ydA5KaW7vl1DDMrr3cfkI8xkNr63nQNj/6+wWi7D+6blGfVJdZ0ssP7rk5eW3X
4+qfgW8BUzYVeM8rslIg+OLG6JeZneuPnaS/tDIClkxKp+JZdy6JOhqnENCSKxgSQefD0P61dXuI
vuH/wxgW7+VFZ9wiwTuvfN3syTfOa8Kv+JyjhwLmAcrU4CBIZf5SK7fy77WorjwS/Gn5XuFWA6Jy
WjbDYLgywX1Zcrog+MU7oh58xgMGjz2VredmrrCKxuzAub1VMZ8QhBDx2S/+4v54BEpNDJyTIqPM
rB5sAO8xUsjYTmuZX2Q6Nzc5WzDkWVD55f9kXlzeGiQfxNy53WaBu75yVN81eJUjjXr99OMAtdgN
+9561ye50JcTqa47dECWyP1RpeE49z90AlYP1EmRA+hlXL0M4Zq39EEZSdq9LMHMHtYn9iFQfzyM
8/aENKcQR9+fw0CjdB89VE0g+3rSqz0T7X+uPhyifZDHeiHqx12LaV2wytZ+ct+Iq/CYl9mgdx7F
tCBXXESEyS2yrw9UbBe8LImeihvi7XrkPkpaPjQwWPiDtj5z+Fwgarf+D/0rBdKrkOJnJMgbc60h
0g9uWuIBRQljkch17fLetkHxlE+hW4mQkHipne3z8H75xZzJXHnOaaP39DEN7KuEoE1Yw6bmBN9k
bPrBc8YBcHSDd1tyTqP0LczDLdJbleEKmrhJWwx3c3e6hXD67YvPTBh6TlD8zSYfMlY1QLDlQVpj
xCPnFqYxIMx/UNaFdAhL3m857UQT3cSfm693nXYFieajACHzzoBOHoiNWx5ruUwFHQatfFrSvu/k
Llkwar57lnf3BzRGCVBwPxJHSoJg6ngG8uHd39ozTpwGDrfo3jDrGtqUKN/rhbncHiULvOMHfsGg
5AIryfI3aDCf+yDeSCPvlB/9JcWB9xLbpRgWgCogjjLxG1G0kGcBtvNwW+supuVeRyGl3n2KicDF
LfbO8XCEwu3ef3xbPKNkgfCOwQBTHqUaYTQvsl4RTlP5r7Zm+hnzx9cAdc1uPdwLzp2ilwww/NkD
2Kx20jm9ycQmgiWxTIkF4CLqIp23nJTfm4/R44Etl0/ZkkpPDzdjUKrQi9zGK81Xdn7utlxsV6Ka
Q8CtJW8fTodiLJslOBR6SPAyahZAtDSz+1tSXqNSPXGf9DBAg/CDYnM4UluHWROUd/l/UFyQZOry
iFE+53DmZOGzsMZQ2MPZGKSuUFpQMIGbfNOVy7jAo8D3CcDK2lx+or9DKUka976//6L0sV0YZxxq
i3pfu1m7osplGXQ9STA51A07WE9BlzIGMe4R5SYfdxJ5Y/bgHiOVCmgmBUDPVDFo9bg13ZTTz0Zs
UkTpA6xlkS12xKwaeSK4OVrBXFClwRELWUVrBhWLBKoEM2QBQIpZKPIuNKW/V/4yiUbd8lft6NuR
XBjEftaSeuHoN6BxIaLlRp3vvuc2YbIRrW5+5sWx3dD46Wr9K1l0kTszytn8w8K1N0BTWyJ+04Ae
eCnXsvjxXu9RVuuhJX4DesOj3O2wBIoOwPQ/e2n1+dUdTyA6hLRDtIZGN+5suFbzLVZlFzky5S67
1vrbm/Jzh5KnrXY0Blzti7A+INNO+1qn+4ID21JbmR2DyMMFDhgh5fhH4vwFdv44W5QPfEayt60+
SZm4xjzeIn45vRJkhPcBXbWQlIEiaJ5w0Zlvjx7gmZl543t7Fhi+CPYXaqtOUwbPF9q5mvAMtitV
5uM3gLVMZ0RB3AFdHJd7qUw/jaJFMvgb2G6tEPhZNyzzk7wZrJlBCdT6gH8YrvEU6T2KZTUka0/4
TZ4qWunrp5B6HRqalsxdHjT5doa3LdNQXZvvMRPBlelwqjmTHFUHS30ofMT47LBthOF27GaIHVuO
pX6W9ZIM6RTNMr+DU3wmEOK69oFgsS7ZGTmHdl+lEiy+03lKHwlNAnv3xAacTmO0bm7qiOmLdMxx
7x+4Jn8qGJ7FGkf3kN5rCbOugMnwZsQZ+6SENMYrd4PoaYHwHIstIFWeFkS41jE9iuTWyXuGFjwy
0mDhHIgULduTtHJVeOhlwKCzK0gsMLUEEErhsk/Col38e/a6xkV5mF6K4QRWgPAf0I0CWzS9rLK+
TxhuTIMavhVxbUF7NMTRCMie1jPEDwuPIEzrSM9hmaLzxfg2SAXGQlr6PgEOs3e5GhOxEpMETKTt
fxEofoX4u+Rs4mOYFQ6GuGLjVYy0X/F7zi4HGF4oJ/1XH7hoI1IDQjSSq0HO1C+Le8NSNesKVnEJ
6ZgTKZFrY1x8fzlclvzMLuJov8rdsCa2DRrRjfzHkI/P3VTXu6Zicw33gBLokZmvvjNria+OR/hK
vXAeUUCzNs4k/StQBGxxNjdayy7G0iR+7mC2/hM87T1q8AHzLzKYr89rGC4+7ozqFERa4BA4+eF4
DBEP5lw7xFDVTO1myI99aQtXf7RR5nfRf5VYwfx99AYOCXzEsPfslBlXFQeArKCELLMC5mU5ki6x
7EWWV2S4tTnW9mpvglim+Ozdg8bnF5DctsBcguHrLvkIu4G130AUmVBhlFyNE2gHGFL+Tb0kBbii
VhwHaLw+iLl9qUS3ZqG57Meg2wiTz87Q+PY7l6uQ2MJY9aZRi0YbzeX6F3P1t0nigpeZBJ44i5ph
pdJ2KHrv23w9xXI8G5EoyvIcloSTqekDM/VmgELs+SUWc6p6dOIHalnKNEn44LDbAzHG629tfVMu
PKnBegH6N7w12F0ubPGC0Ei3G7CP7x/6MWhzS22tjTFl57hFW97cFcTpj+o690qdSbVLzHu9jhYC
4d4vDrkW6WpX6GCA6Xlwp7vpzQUiCWLnbztFL06PEQnYTbKI+xTRLnego8L/qtIGL8TM/wimeYyL
aOazQtX6TaO6W8IW95HgpG+Xo1NF8CcM9FDZ9Ys2qe4HetJMeBjHnGNAbB7QSDMfr/dduy7KtngZ
c9MyEjcqdEYSskNI2C6bkhqWV7z8qQumNQzENCWgo+cM05ybkbNbWZKdaegd1ukLgS6jvKeDdl5v
H48QytSElVlkts/GQNunIk2ustZCCuyDsr56BFxf6g9Ut8yOB5mr6CfQ1p/WhstfJ/pxO1WIFE5a
OXwIrCbMZKIBqoawYGG8M605m+55UmuxykJ/ODTauKeTTIUP2YlTTZNOFs2KomXIRkXCtPX1e5ot
slfBcfxXYSWSX6sjI2oHjMKY4P0ejX/Sk9iDG21Js8bkKdLO07wljSIOOAkV6RPj33TcGzVs6RA7
ZZRVQ2dXhoj6LzOa7TbSxFweMnNwTIJF0vR9fSKk9Do04qOkM6cxn3N0AbSsAZXBmhrwMUuX8uwX
GiDMt2Gxo0Um7GlYESn7SCreD53uqCO1KJUGjpxeN8OjfUzaWxWVHt7x8CaLCBBlhnOpSFp1Dm5r
kAFfa62qHL7+ybJaSa5fGWkEB+dSrCCSEeCnAZNjIT0i2goA1lGt1yyb76QZ1fLEEoPgT4sceHH6
tycFyEpUDaDEVy0R/keof6X+7jV3FkSW6JKzWmcvnsqt89XLPV/4xF5nv6bcK6fAcjth1VvOHHfF
LPdHriSIP6/lUVLsMK6pjJl7HxV+eutKWv7O9HUDgg9M0CjRlyz6qAiHPKb8sXmOCtYR6F9P/MqD
9vb2IBE7pB8UswXW3K7L6c0l/XJmYcpljPzPU6hHNMna3VQ96QD1ioYU5/IQEdAxXV7mOSipSWS8
KxJVK8mhxaiQrnbQNbjs2gdJrHIRvXluPnNxZqjPIRO4C7bc0+p4iaGImEViVEZEexgb0CcVFjrw
h2E428JXaZWNKyKV+E+FCKl+C25nwsrrqcKx1f52TxVJlFOkg6wxs22rWwYwkM67fOEbCSNJpJbw
v4J7Fx35Llpw70YuDQ1ZqB8H//nSfNlMR/ONTwKUd920Tg6YOE56nuv0H8K2kyl00xrgDlzuTi82
miSzEuJVokTWe3OSSpKwIy8QRoVBx9mYahoQRieRYNrBeVCxCqD8ATmjbgXFOy167nDudoDmPKQu
qNK4Niran0cCtJ4TcNKnC7VvqfRHOAW54cs2trNkOOzEeUyXabmWPZbwcvjCqCFYRO9kBKZSGXcE
/upAZC1tgbSmuxlp/3A2rhZnyyAAXcagQf2a/vvFoF+r4dafCug13wlGbEyondPnd0y389LDyn06
DSJocz2YhjFt0hq3nkaYgqeon6BwB7xy2Wd3FzmiWs4nrMq34CzpyseOLUeoehGZONHFWG8SHEef
gIBXSI8Cw8h8oESBkTQjKPbFGtcKlE0GuQ36VLZ1wiME8vwZUsBpgjJ4Iu83/ar7tSysZqQmUUlu
pjUhBtWtL6wt/MYx08AhV9UvlvrCFFVM9GEeP/OPOkYPxkRGLPO/Ek8jiSlfRwLupajrFes/iHKJ
/joqVMGw8jYYVjhGPsmD8xld0jY0JE+oBMD+5KBqLhGKgDNS4/nO9TcuaqDCmzwcthBKIjyXEHBY
C/1/8ErUDyO1SjsGx9/Cx4VpxR6ypHPB9XyXf2GAHhH7nUFZP0RCwSeaUGseTIACtUsL4r4TKpQF
f2GjEeQd8BdXMQELK7TJB0X9E8/R9bPOVWZj0MjvQCgB6+cwGlZdCParKY66UKn8jFbuCvDR7jfM
17jOORNhHX9LCBL2mfq8KN1/1NFlU3HXha+qcYPFHB8oij6Fecw+R842WPXdKyhhB+8/t23v8CFg
xujuEwKWiSl6sP1oY+HyV+aXeWlLlaTOLb+dy1iz6Gagmav8ZTyGuMGbYwBjaWv6OkOHpJYOFtpp
X+SEbCOaaQWYCGCFrkOFREAI6Uzors8aG+JsBJdsAKYG0bvhJ6vv43yfCul3z9doPOsc0OaDI6Iw
+9a0ecU/wbnONx8m1dPp8so4+wIQWBj3Yde/SZ4PjJEUTfhsV8UZ6UhkQB/AzUaxWh3RuFT0WIPg
x70RKHeSbInqDMAiXPxwlpCXQAAgVejUjOGXRiQ211gpgyqQCU2ughh6byyH3Enil5eUZXaH6qQi
sE2e1asCevt5gdd+SSNK2hIrHFMZGX18jsdDHDSie6IzeQsfzuDL4tHJauhIObgw+1VCYAX1gEjw
g45hKdJtdWMBFUUnykwnSvk6NlxgCmne0UJaAle69kCWb6BV9X5Ple+YLR42UK+WBDLBun2THQYv
2e9oe2IWeVNbepHY6PAqxFjScW/Uh0viNP7cJSbX9mWscO/nXIdgto0aZMKLp5DYsqq5uoSyd7fC
JGC0b+fqtmjDPLCOwZngA2h6ILUotM+RGj6ZPG9U1HS/OlT9gFuNcLZTaT0mxRCnJyg8szC+0t4h
tWS9Q4PkaaV2G1h++Y5UWNwY58grX1fefeapQ7D7VlTWuVpj9bTSUxm2fyvo785XywFTo3BycqbJ
jMSsskBHHBJ3v7h+WI7EcK33AmJ4LjDN+E4GrvEIXABpkFAkya5Z04gXQpJEGh1JP44brXaQrUtY
I0OfXyOFtsiUX/cTpWYoxJGNAOYSTY6mI9sEIMlY8rbNscTIbrfi6SiGP71gFsPQNltDpRHfHRuS
vcjAFRFImXQ1rN/zI2edAE7gpcwYwixchp9h4/CfLQeZ1uomNHt8jZq9CppZxmsIvD47pkhbpBB1
BgGZMI8MYtAJEpz+7vnvQKAAxP6pqfJpw7oyL+fwhn1mh380nsAJXV5ygi80eC9p5KMXqV4mD8to
9+1EaYSoNrqYbm/YbiLzkzuxI7dkz0MJJayeo3JfA+Xq5Aj0LCasfREk9ixFLZYSn/hqReF/c5W9
JBCkN+4S01ruCBF1FRHdoSJU58+CHmxPQQRCuM9Sz/+dHmHgjrZMUFQkmsBfuCdOIjghLcUN8jC1
T+pxMlnrSGIgods5XbtkmcatwfG1svnE1nG2qsQPWUcZ5dw9kPvotm0ndHNr45k69AuOpfTvBo70
OfI53CnEx+TAQNM+hTEounEcYRCg3dl7HxAn83kMBA5xPw3821+8uI6pAVahh1eulIVoMQHKiOfb
Cy/8wVYnEjBNI/QjU/pv/vV4lqEuIR8ks0KDLOTfOTzLGFvy7e4MjGmJOYsfnkRuacajTEp73Lse
AKhzjmeeMB5q3Cjmpr0WW769Px2mOqoqrvNgKRKcrObjF/pHuWFV18AsvzKEyDWajR6GDqC5qGRO
+LdzwqouIzxbwN17uhGRiUxNbJ06IcbOVF6ZIaxy+6alGDvCUv00CnB2zQpnk0tuQ0/So0NgWA4Y
owyqp6K6rlUcvNS4tWyX03D/QVlhsccNKSqhwGXJofq6vY9P0h9/BX8PK3qZZTM6ymP52vIKeIGD
tLdWT3SnsSl3zm4/LyTIHmh6iB8CcGbzqKOhoJeTrr+SkrG4E0mqJgp+4uHtSkUek7q0mPtUV1Mg
BBNoSyVfC8Y/cVW6QQyPCKkKXNENDI256NuPtNzj1WCPRhYtN+xT54F2gQYN0hfrQMTkgkUGbofi
cTxrLj5TuiWXbVqfLa+IiyhAkZZZngCi8jq9FSEzDWPRXbxuKnJIJuLu00hIcwnym/0/wYYE5RyI
duNThQaG4iN6yMnuBFwgwHLieoDAl3x1hEDWgzNylKBXBeDx2wnQFTZit0Avn+NvTjHvQEhM4PKf
chC1G5d+Hejb13XqGrY0Dm/6gTi9abaS+hqhEgq45P6yMzB+Qe4xUEKzr1Sp/PUDUa67ipEtCFJn
3kNmbomhxKDRlVjTcS8isU4CNfjq53TZ95yWEziNMGIPrFtuRS1qUXSq0ryNDqKWvxOoJtzHbWZ3
P9NQrA4mXidz9TM1DUnvxH4L2uu3S/tiogQcLKXFCVlyZ1GzzqpaFxtCg7bOdzmbMocuAm9O7Dzw
MEQXt2ICS88jAjIQUJZrm6X/PkazTij8DFsy5FWEmI9zs468KJByJM+tjLR0288265/IZ3ymCArQ
VM8aXMXyp/cuemtDuMB2+9jr/3P41ch99lYdWt/yk4lofYujpL0sCz+iKs9EpgEJFEBQ0CcSQzXD
uq0ffYSj1D1fCxt+YQOodtxEh7E0fHV12AgbbcPi/h51emMQWIzwnkoG+bdwq2SzHRmdORrGQCGl
HQXvHbdAIBAQNciXEZtPH7U7+ZUe29WkmSHi1ccYZAypgxrbpk7R5KSq2y12RzGZ4EToJl87JRW5
oqTxUydQ8MOD5II+RF5qijzTtUhU3UFPoU9IOxtiMeFxOVWvM3YZT+BloQ7s/QacewdNF4AVXzxZ
kSPFqJ7eA984uFuuxFepADk43o08/R+cqV6jdEClJXXJ2Kj07W+nUneUBg8FqVJhbG3yRUW20gLQ
mw/zGVgmlTudCl1lKAPa4LqCoKdjK+Q3tUiheFAGUF9cgVj9E9FwVd93rusOobMSXnkYGqYZd5A6
E+VTztXNJ4KpAEJWfLp/jCyJzgD1JQWWDrhJUF6JLHjDpdSd1xbKZJoaEu7gkYpMdFdsn7uA6Fzb
9/ix5AdYfNlKnMEkWryk0K0dmJScyjJLD/dVZWZ9tHDMemNtj+9p6iOG5AdaEbzbDXXVisuZ+w3J
d8ZIHT1w8n4hdyksZXlboI1ZEZG2+ZRqodmMxBogxxKbh9CHwy/vB+nS14Jjrf14m5xU1Zoqixp/
0cIa0CWS1+eoNmV7PPWlJHhMyvMMArGDDLH1Sk3tq373F3huZLz9SR3xSWYkxiemQsTaEvczVP9i
tTV9m8JMAAjJTWmGdxqprpK0w9SPqlyZX1MPo9PM2jBSL7Fa5Qz8ps8dYIoW4pb78Ws32y4muCxT
hPLSf8TWQ5hr6MAM3xAJ0ofdnC8Lu4x9JZ/jw+Xk/gJzNee1NbXMRLfBAprNjGg40WWNc804i27B
ZbWaD1aj8OMjXRE6Kah4Z1Rx6IWRQlVgBHjTnB2BqQU4sTenlODM0pncGvRjg/0OITQC7vG50+oD
GGVhS0N9Oqmz0cj2IKNSu0OImhR0Krc4n0hVT0rZOsTUAj8HCVp5flvScMqOZ1g3+QDJMCLHMYxX
nB/6HK/m/KkuImygKGsphcsPcJT2cLDGClmRziFskOglfx9Zys77jnWUcxLDhPOIvTqXRAV6CVU9
YsKP4Nf+od+l+dE8Qb3yhKL721VeGoSZ22fvHacZ3Hqly2sKuZCRxfMawmoEztEbymnVhmx62lr+
bETclIgpILm0ZJ9+C7xlPfT+M7vESaagMWwBZgLBc/yUnwSgyVsD8twu1LiURVxo0MfdwzjJT8JI
RQlP+ygB+spakYzsoN73F1QL7VXF69oVYNNF20tiUoTOoUz4WBtWjhXQ/79oqQHn1Vbf2pvjxtl3
cRp4/mbsBHIgTnsunE0aApvro9trXQCj6E0NIFU1vVtztbUBfnXTQ1qG4EAp0KrGqB+OxshcETfn
hXiuASQAeh4HhReJaTObc13Sc78qOdnKsHp0qZ0xyYN9zfaJrcKi3+3qN6DcGLrouq85rUcinOVz
P+3QGpJt6+chhKYDRm1xjCT3ALhbAfZPx12LaGoF/NwkP/Ke0jGwpTP7klqSjhqkZhjkrLdIS95y
MDq4or74Oiunnt+XV+hX20E/lLZGyMCftTLXk44ctqnugTZINWGU24tOcaSoXXwj2KJj37CA03ec
fV3hPLDXTmvNa0vw3WzCY1FP2bmcUZT33U3MfhNnlYQM90RwJ+eJXolL6JM9fJpBAc+u+KPRKs/3
1sd1Xj6QmSFuaftKrk0sjqg1vaNmQc/tYlg4VSBDfc8fCwWqAy2CHle5L66mMMGZdlj1D5i9KPWN
iVsyGSc15E2SAoMVS2/iZquO2R8OOrrAElUOSh0lShE18kFg05CSKic1o0/X0B/i8TQiBg9/A5PE
n/p2kTV0lJIZLKhZAkiZyDTWuSnDYyLxD6+4Dpzhi0uFDR9T5CFTqxTjhB52FUX4fRlLatZ1KC9j
sZmOPyYG90aVrjnga58OtmPO5atMqutzI1wIfAdyXv2iLDn6cWCyB/go60CQgbkKhrftgkDIMQsW
5HI///gh5h9nyX24BOZ5YzxvGDDsOyCSGAsROEc4zbGpcX0ZiQnQR145K/cwIaZddt6iE0rZfQyf
rSodYKODbsEAV9BMkhIrtSnXDHAknFvKOAOTT1b986PssNG53CtpfAgKmSTosoPx8W4Bnj2/GzqX
v4xNM6a7GXKtnn6HBVcGgfKgOWLq6r+f4BIL+IbuUCVq7XxiJ9fnZBdhOupsCzVLikOLcGl8mtJE
AoyL1VWipQkMHdhU1WEn0VD5mnloCvXnOAeZJGqUECYNepIBkvLxLDEDLSndCmD6ydLLtYNF/9Yg
o22NKFRkUM/8W/DgBSxyon7HtzOX1KWiXRC6iS/QAs8Teeg1SMVXLJl0GB7vr4g3j3Dbejd6ANwq
qWMK9oOLHyAzC/cYHt3ZogTKkzqK3axi8E3PCTmGofaGmj05wXKWKJXe4D1tbz0JpwzjFAi+NxV4
Ky2wLfy1JwDyQ0yrodI0UmOgie1NXWi6sw83zaYa/7Y1FNceoke+KIm8D5FXpu2NCE6mYA/m8Cuh
INTQ6r9fqYbyq9mmUdu/BQRDCsaHbdstbPfeKV/1KR1u489GaYpu7rMxXem/3OIfJ+fZs0NPKjW9
bBu7BAaTjtayWTRbzluwEOoGv4X8yaFSBmmlQbtkJfCkTR7+K57ldk8oSGjeKOewVurEZrMCBIMu
Um6WZwMoY1c/z16InTZ6ExvKcE2mJwCZl+GkwwR0B8uON2K0oteQQ+jAka6uEQfiLQacU+vEDbQZ
idDyKDbTbmcBypc9+65vycTkYl+tkBmTlrjH6MCDL7sBWiPl8OaExlSDwaw2UNCdJ7eKWug9ZIaA
3LE7pWY0eqxYEWmziTRF+JOpmtCDXQnaFuXu6dL5s+n90OkyrvalcgEAX9qCUO3qsvXOlBS8XF+4
ieMokI6qyncmTbc4vOR6SFRkbUGo3qmimEuuUh30zrCbn49Cs3OBMPQfu2GATP1dHoncQHVroS3H
R8dNHmA2uKQOeQB76AwJHtNj2fnMcsY2SH2Rj6YuwSipLz3PUjgy2uP19fDsU+I4fiGLlSDHp2N4
OHSRSkCVjVCwcKt3LZEZzeOIGFc7Yim+okV50M84HIpDKLUIqXvDL42Sdrz3+oguA1PYhSlP800c
J+6EC1KgdCiQRUd4XtrXEHw0NAhZZmlWFMZPn9L4OOeslFSeBUKtJcE/NEIBPSMwlIvrlOrkdIw/
XmoR/x7WxevVHroXxmO7tb4zG/nBJdayp4BG4QD15079xQ2YzmvsoWAZE3wAlJR4ANT2M20WtLYG
9ympC5tJ0ruylyhWLh41PX+2RVhBf1Wh5fFeLmcNPLZGS3gUqA8WH8ENyH7V3lLl0KH88Qj314Z9
PalWE6AljiW2R/VQsBKoKbr/fcu2YSABDmGNkcDOdrLh+6CbCeg2xGNPr3pGDymKfnJ5eECsrIXj
KpnoO5Sn46WvlZM7B69OxpVF8pnPpJzLDwiHiFHv6TRjD/uib1nxnV8JqPS+lAyO5rZNi37Z+TkB
C6P5SUAZFThChpX6UUpKuYip7Ecuo94YCqgaAfgDTzgu4GIsZ+lRnet98y5rEo7ISgkpVC/EMNZl
5duaLaey+u5EZgopI4PGTL49VgqxXtjQfuMnq556qv/6cHJUB98JnRbW1f7STJZIS/8entnLJ0JK
nndReXbRREtOKNYuUWtsqNkDQH6Px8GmE4xc1QLDZ0Xe/GMt3wsEPa4w4dHJ5TGSyCcHgruDK1hE
Q7hn4XQYS9HiWkYJmIv5IdtNIRJRvFNkcd1FTIoE5VdPV21cQe3Keb5ubw1e5O9gppnRDW7M3MUq
r6EwQjXBs+ycbYEOtZxdrV2Y6bK7RG+pntg18qQ+MB5zfMknAs5Hx/yZzLkPoFiILViAuW3zSvHB
vkbKfrFKVLxEtS59DAemwkcJo0as9+DCOqw29wDVkzgC1TFmhvC/4vivMqW0XQVNMPL0QBiBa1YB
ChZz9depe8o/fwDTAsHDAY2MLTqIMCBCzHapTxsB40IDOa6/o2225rLwbJrNzmdfBDfQTze1CcV4
qtQhij+h6MWe2TSNemNmfcaCC1x3zxtOpCfT4he/zSVR0dC1RAkUV4EUUBQDO0MR4yFewZEOSxta
fr2ZRls2jTQDd8zqJxRNJoakbuLMHaoBHUWbkMo9Q8cCav1y02r64QMUSM8HVbLzhz6GDGQ/dhlZ
qXYszj3qTgpatYh2GM+vPrjq/qM3RqGDHzXqx/L/9oB03uqRVlW1FTfelvWIqRKpDVIhJZzOpxV7
oytWHrzop73lyyaKw4iv/fjVIlk2uTKnDCGzZsHknFwzmfGGa6nS/2+/wHohaFvJlr9OKURSvLDA
AsuJG3CdjzO4j83Jc1zHj2KzbWfQ7BrEQus0gi6VFhYanmBUVOVaYT0FE1vaD0Q9BbBXsBKhMmRx
m1Ko6NVp1sdrXT/aOej4C5Fj/NDeWwzq8nimmXtPdwdTUaX2tFZMoTSurSkkEpKwuHfV1f6SO18F
nkC0npRNBefrj5Oilq5ZW5+Wr1f9r4pEJiY6G9wWJ3VoQU/TL66hxSeY/mEfCqxXDPC94Sctq+Qz
5ew4Q8WCPhLWF1X+kt8qAuVyd07SDXOB9X2AdXt6yzL+uMphz+GZsfN8NhPmE3meHOpVRbrxg+15
cUhAJHqQJCj0WG1pQ7xnhYv7Ujj4F3bx1N6Wu2iwt91kzPWPuwzxfg7AW6TCNP94cWFbfgEc43xw
L9epObmz1+hDWVYJtl4Zc2gtUePHc4EwKWoDR+p404LK8Upa0FPz/EwKjwUYPzMC3U5L4DU8Bh+2
H2HZpF6DRukk79faDq6ZZWK6ty+52N44AYlg9RxCBCBwASm7vAtkQjmOkaGCTEsnPGN5j32pClPa
LR49ipzPZuULQTKxI5DT3r/JYxETLZpH9B9hRfvwDb6LtoTTguqSbB0v/0IFCOe492oFuCVhgvOu
LAWay4Oc8ys7bNQpgKOpo0B8Uh1EogB5XqEz3T/ejYrhnxJULUtDErz2aFATZYOm9tKXzl05cOrI
szT7HjfpPikocVq4MExupOrg0e6H34ZMQecFqarimYt5PwKZ5qumnmPgS5FcWjVzfzVHe3YR6yE2
9zpHLBLxgttYnThDr0+zn/kYN7c0vpTXedFFr6fCe4FB8u0NFrzo5UvlNdlB0QcpPRj2TrT3mcIz
S3YtPpItj6HjUHOMK1s2UWgSgj+Mp3rqxX38pEKbdTQvaJQNT0FsggsxKekHA3qSmcLknWNoDtem
lkiAn/E7zpmwfn8pClETV393XA7gfM5L4jxx2heMYj+ldoWqyKPt6qS8qZHYoq1kvhD0vMNkfTW4
TUqkSefZjendO+NZ92PksjzacblfYCHX0yR76HHSv9YEuRXgNwJdGEXSKCTEbrnP3y6XzT2J8A50
GZWyq5eGUuGQOWpBtOGmTP1tgAA9G2HRy6qvX2GtX38pG61aFRIDWxeB8Pw2323bluftjPxxOe5O
MRPGChu6BuFEInOCvBfZ/F843Z0IBn4ZGXoIl3dwqKPC8zt+qHP8FitalS9nN2OuZJsw58gm362v
KTTeRSr2YFfICP7+fj6cwHk5iFxF90ViHgJZS8Jio3YHdCwLLeJ1dPCVeEnEFEFIYDx9Q5YoYNF0
laoEa3m15/ImSrqJsVs3Xh4y6OP/Dl4O+4heoQlYzKe4ze5xad9bVhQAy7W7QhlZYEVropYJVHQ8
EgojDdCYUigtSykkVA583b0YAOechJ8wyB+uibOXEnixFNy63D+GiqD/AlvqfMb1gfcbHZqbe2/p
bZxqGStgtFPC75dsxn9b71nN4B2xz95AZT9f6hZmomzE6WdIQ2kWabp+mpDDCvI9EGV9zvqzxRro
Z+QDx00m0dvUlVox7f36/d2nTAMey7Fmz3i44tv5xHyNyskgF8Es4IHhaDaSCyQXhlbuf7QycJgP
lrWCuM8u3ht2PcbTiFrIwNjJ56oboujEIH3h1Xb6fx9WgA6t6PyZzu6mFZ+lt1VkWlRStSRaew4Z
xMuDBkQaoolXQu5PoFUVjgsLaNWbehHuw+fcpwIHOhYbS8Jmzf77UOlRHjZfvB+DAyIa/J9A18Il
YPGyvu81mB5yFQwYrKz8twGT0sGY4PAKTjNH+wzk1J02yV4EdPOYlLaI1wNF6QyfhbwnX6SKLs/a
b7X64uMysFbM2I0ojc8hdbV37Jcwro/9+ilM/XIOac1xEzH4X5QtI54O3c4Q9UBHeQQNfyM31Kd1
P9KDfhez9NdtZ2t0r4SKemMhtxNX9sk6HXMMSEApM/OaEXQrKpDwTFl0Kt53wP17sy7mqByu3N9l
vHLWYP4/yCxImOuqiRSoLBsmsiMYpmss4KkXn0xGvEabY6tLEtk7rOBo4qhEA21948S+NKa/kPiU
rC7kUPENnH+8k45jCpkS4ZnxwGJGxGcs7erexamRvHge13ee5RQmL79C5XZ1f9wx9/l2jbIPWVYX
s7ByA6wG+q2FOLeYwiAui2+tBHzLBTyRzbt7W4+pSLpCEnKkPFP+QO5z9l26UKN2MlJbazNvWh6c
RH1P7FNtNpgkP25qyWqyE39PMe2HKvxe8/Kjy9xRJDOj9NElk9NhIx64gb7VO0VmpzDGaAbarGUF
l2KLYNDWd9sHuHLEUY044lMM5D9zMwCuV5EJ+lDpQMtJNfqYi6+gqyk8xyMpxvLMHIZ9dJzUUcrH
GJ3nCkHW/LkZMGG1pkYkUXB/RzJPtw+E44DARIses/5xya11754aTJJR+Q538GDiwNs8AuvG2In5
GQfgUr+CfDpG8PG4ZHDpV0pTA7pGay7H0Mb9lqmXCkJQM7MD20tDpEwBy2X8oAoJniAJYy1pXBmC
Da08PG1BB87TAJSIy1V6sV5+i4hrqQ2nUFw9mbvdEj0mRCHczdQ1w9kZtkwScoishu9IlsEeUHCo
1RmOej2qOtSiX46l36ccVe93GvG+HlsFWCS5MFEz9Ebr9j0PS6RDtv2GyJrlnVqlUwu5NThjoqMU
OMfqheqJAVr2hc8xRQQiGcIINP1UGMRCpaRhfCKO+wwcmIsrPNpUQIfyQh6u+r8FlrAfskNYLQ8u
adkr31DkTsg+QBwRZwsN2imS2HtzTOD2Db/6zbJ3b5mDdtjAfOQ/LhlVHzry23/Ry0fXBumVQXTj
QzqObspUIUtAmMp86Utsmkf4JMHkJZmaJupM5hgoqzys3TEaw0NTxRXr223KXzZsseoND5b4TCHZ
5knLc1OFahmj02M+lcZJ0a81dsOacP3DB7LQPfG4POw64n9XYR3l3pYb5ijuZIicOwceR+iL03i4
O7YCKYIA2CXZQA72m8+v4mguGeqyCu3lh6ASBhDGlMSFLd/qbfMh6aLPQCH/5lihOAte9q34r5EG
jlJzWX8UsGOhOdIIo7FziF5asgdWpkKCMV7ssA3D6a0cdrptN5e+/18Jgd0ATU7HY7mtC9Q+f5oO
1affTkEV7CDZrKbwIL3N6nvrStmoRsrXBJJsoxd1+Z4hdN68M/F8k5v9gXDU8FWwZTqxA+WmzlAr
sMNsvAFm54iqIGjW0Ko1joGvABNyRVhXYX+fux3V7xJKCnAmqR2Pch/Caix3HB7VCnNinlskzBHU
Lx0Hw+6SOwyO0IHOjfk0f7GfuIgm2wjr6xmqNtx0rZM4MN8nW6hzzJdPWeSuDQMFTs2F7Q1JF3Hu
GYk26JAfekOxNKpM7hhAH9SG5RcjDxD66tEA6IQcU6iapXO0W++JkdSYQQTt9JSH9BxEqhdgC8JV
DptVJpeieYoe0t7ByTH2g7n6nufSn76DO8ZLNIrDkwn9cdVqnGvOiqgsoVg/u8p0x9ow4Sct2u/g
D/PSUGF5A1mgwQrATEm/Oh4RDtzBFDUIZ4AtFtdiU3DfU/DUMfoX293v4UXKev0/HpEeXEg8RdCy
DaAyE/YRRAT6HHeZ55DGJDTGdaDmvu7qGhmrMI/+scTAs2ga763kZWKc+BNvZ/oihj2MicuXLjQu
BqWXDvvG24iTt59oL0g+Gbuwp9IPBD7PwcBzMjaVSSFr+ajXLXTE+1kXdL8Wwy8q9xJBRjjE8cnh
dh1JosJcq29cFswrsik2WT2OXc3FWKKrfOPZF1qHwEXWK5pGhN6Vte1NvB1Zo5zNm6VGYBvf0NTe
nrOvK2lN8ZU/xSIx99x0b3hOgm2r8mu2kab3ijwbMKTVlkKfiWTXcYNeNik2zoXUTcjTtyDRwV2z
DoJtuvlL259r5W+kWcmDtlwVyJMkrVCfqoXVvXwetp/q6DqLiC8fKfuqB9OKhQ3lsJs9X60PYMzz
94iV9B6d93Kf6kHflBgXsjLTTSzXFM0nSkCI3bqrh80SO/y5vSlhkTL7q1oHoV5Iqlp+MJK95A5V
qz8KwZoAJLVXECuDL5nBDgTrIPfPpVBtJOtk9ICpRyfbEUSaivVQwS/sHB+xal9+BMsQvrlOZRzf
8ZPZYThCTaKXHHiGlM2MFuFkRqZs7fRPmLQgFpYLZ8l1Pmokob4Lk2DuNih1HiEQHQycmo2kpjhO
UODVonc9XPYPM4HsCtL4ibTC/1wv8ZWpjAG9EEWGximbI1tvhUcu1CykYruIgoD4YFygGhVi608B
dLuTuq8HANdfxWcimQUd7sBJ2EUvy7qHqCh5m+btws7MyrjbZUVXEw8GUlwFPWkS4PwigWr2J0Xt
sOtUm+t+XIwEIZYAM/6bAvujSOwJxHWKyWcEo2vrRXPoKL3DYShGm2BLTiucBulMBiqzSI7YjnWZ
iGdx6IuHlnqAu1KKM85sneZiMlHKdmqSFJ9+tTtLeNz+/KQY2xvAnD6s59aXxEmMNgpNt/Wi6ewt
+YRaj9ujWOIoA3s4Hrbyrd+2ckARFvvZ8Qd81YS1R3eUheoTkv9aX+wvHDSKm7f/UbPV9OMnGc2J
Ameai4WgpvwJquZQkf+SkbYcxh/JqLJjotiz1Mm7xr7OdZKRf6ZsGsIWf7bt2e9EJnPSNcSHcGa7
x2JV8uM4FL3hfEoHwU9byKIfvh/qRoxalmP6elJy+KcF4w6Fx9Ea01OFK9VN6h6MpLMo953tytiW
1kPfaE96Cgp2DSZDat/evfXueoc9aXC58n2YgBb5Q0V22mNxFk9MjWsoUVOiS/cgRrP+SIVZMtKf
yY6HZT6GDqF5brvTfYk30JRLBy7omjxPGJlEHJLsQkQ/sySg+bv0CtLKb2dLvA+W43jS+r1FYL3x
+vhMexq7KsxZT82u4REjrFjYyA3OzwQQo2t3sNzrCkdZ8i9wMd5hKZjuIaWHLFMdRtKUOS/QDZlN
p5IZeMZfaMYVOqG3DZUat+ZgqgErpAt0LVrIbJNFfYMlkMt9cl9GMl8SRoeN8rWn/w8gfd8wo68P
9zCfhDwqlGprz1/F0Oz6tO+NV3pvFeLnqYDsKIfxCElJps6Zz2U+DxzuFABHtijx72VyBKzOLb/4
zaHbhkbXlZkNDt+YyfLtdnvAEUCc+x/ffWTS0oFW5sFSrxIyPms5pnhGULXyM8hHUqSK6FG3woec
B4jYDnzRbYnKN3FPZl9e0UHCAHhVl4bdPrwKCCgRtJ+ZO2IE7VbhHkeHK0ka7OkCE145+O7TfM9H
JjZ007Gm1M9D47HpWhnpfiemH6fwgWQzsfehuGr7//WVak/wJJVFiNLohE8k38K5n9JROyPFYU/j
K01ZCKpi4VNQg8KvrfLZXzY94T+j4612bPqaYFrd7fgubIMgksuTf14R9wUN+Sd7+fwV29lK8zmh
Oeh5A4HpIa7KIwf/7nNlUTgITo+dKFof2PHsCBRx7+PidpJ4BSxk5weVfNNDm2brBPtwE4Gou4Kn
DmgdHrntsDWx1w2EKk23KGGom4j3SgFVvHa+LD/MZJOXR3kIfmS4AlZCCQ2RM4cvwftRkDXuHAB/
vJmdaqxQVNrUunaw7fLjlbcKUsI8GtDynHJDMr7dvAhcjUKG3F0R0FZt2Sj7OTeRnjSYXQGhcOD3
Tlmq6V5XsiLXQj5d9xpSz3W944j9RvJwlzM3MNQW/kQ4wuhXRz8fg60Iok4CaMjbmARpWldAl0mD
RFTh4b5P3/WDHln7MJwFZCp7b+yNjqXc5zN+ZEjmlui3C+gvvMvW8Sp+PamBw3HEhIYdPsl3i1Xh
R2nAzYR8zpdCdRVpjJTDmBYfE9rENxROeMHlNt1KRQcSfdrZk4MfJhzrXwr9tIo+tQOABGHdkfe8
K51Qo6N50Ypdf3a9VfyzmO7UPkLcKbeHa4MMX0b6OF73b09blQfGOtyIg+XJiXITSCFGL7DEAACC
vC11HZT0Ny6sQSRFBXQSNsS2Rrp9EYqkqtA/Ue3VJ+Gbp7w4oNjmHF2ZHCb+Lkd7vJNT8T6NF7Mm
XOyY19EEoAUW5etKZjTkfQXzfE1A0MOMOYdcUtdRyTYFKOP9+rsKg3slE1Vk2knbvf4so4R4ZTEe
hE5By8iIaeY9Ewr/xPY0AtSZ1mXGpWXnHo1L+Ak6I7QExcPNbPeR0+Msyh7VoF68zVmHo+ab7j8D
yhUYwSwOdqCChjkCjUi+Bv6AUQqPjRomEghR/C3uJvbbZWK2hLbVXrKyTqXKZ5Qf4FR/MUu8eXOM
Fstv4+z239IN3qDoMnH+Cd8bItskT7lQsLk3RPTPbaS6imQ/xClybLsPk0XpBg8S9O/8EQp+EyMA
BS+ZroGsZJpmQyCDMhjbSJdGX+YYrxzq9SBQ0TdgIdXd7e9mrEVhlg+KJj/ex8RcABXDEupNLXhn
Poni7RHko8as6Sh+Ne1fQRFNH4ow3LQ5CjED7/p7iMHuqeLxZjofYwofukNyqHQm3qYvO8+mQizA
6Z/FHUcB+Mye8Ex/tPJeN5fY4E5lgiD1Vv+khJDf516T6tjxs3Y4C/ytbWyqUBVsuprF4yVHVrD/
yW7kU5sMs3iYStmCrKdzwuzbBFLO7tuaJxsmXh17EQCSliqIpq8KdcCtZAA/0KVqPyH2out6eZ51
/3VXLYCoGYoZw/9IGqaTQDJfKu6OY4QVa8ELNofTbIkM7lar/nnlXvrplajs6FB0MRA/3ePDczEA
Eph+X9K2tsk/PXfxciuCw1EkuSl7gdjTEjTz6rywU1pN1ZJ0IjCWhhD/m1ZOx/QFRUeaUCfCARvs
GWpi/jYYixH3aZVDNjyiuikIP3KeGjgXfTXZ/2+PeVGujEcLBqz3sRKFqBUPiawy2MXZkcApoTG7
Dq/tpIA9kb5TJXDRE2fmavCdbFfvpWMzeXiAEy2mEoQatN1vbHSYD1WnWOuNyemgqojuwtf4U3/l
Etk1I/R6wjgR5LAHd5EYAPQgM+uoV11sziI1IBU+Aos9uZSpxg4oKRoXMHJDITKVBucMHOcRioDn
ZmwhHV+7ovs9qsUX58B3UbwWQPiprPkxPBZqEV/BxKSgsN/Y7Mi5ydp1R1jcXmF2c7HAJy5ebnDT
3VnYhAt9aZJqlOdE+psvvgTXlW9G4TNcXyDnB3SOYl3aIDz5aKlVuPE0Ug1OOFnNn55MatzlWaA1
AVFPU12+yjrqVM/t/UfnyU5na1LIFXnERosTqlK21egpOM6SRcAmpr8GtnSlRdLg7jF//iAlo4ca
MpNHYme/6NA2nT3eRpZZI1FBEi1UMCYzozKdF4h/sKQD1E8bEzdQ+upG3qoI3C/GrYnaEuyRt/tX
BXtTvNBHf+TF3QRdkLitA3LQI+9zJKpWP5PEd1i8S7BgHyw/OMjx4iz+Dr2si+swbcEt0wZP27Px
jSVFehuIrxW28rZGBX/MAUg6bY1C0NpjGyHIQuVwUVXxOCYogkUxu5Zw/QcrXzwiMrKWDB7n8W07
eBeb0hBX7U0zibBdbXmlL961mcYHBMgKECxVWxwvRUyfy7DUGHSAck+NQ7EViwjM2dhencPYsGSQ
+mCPec3VkXHkmV7rvR84bLsQqv88wHhX5E4FZD8UJweHhJ1lI4itvIxxZehJwdlFgJCd1gxzrE3A
px1Osem/zid3kn1SzFaHfACWjdjpBqM2vRQCwKRFzyySajEXvi3Bhp8XGOE8SutEFE1oWCbkoLqV
Au8c/IQl9YPdEKG8rleOXX9M8lt1RzZS0XwC1ekHuniN6DNV6sHGm3GoaqMagyUfRYgEzz3ieQgA
3nQfDfraSQ04Aftjf9Z68oqeww8axdXduRJPv/o20muvz8KRtCqTPMBNZUBqiw+d/wnb6bxrNL+p
6lOx8s0+HyofPwraAC9YwGn3vBZnOYRlurVmCrLj8TswmmTWKi7LiX0zzDyyKxFbKxB7bTBpvCax
FiSBxDRRA2Mh9K6E1UyfkD7dv82y62tn+pNnGL5fpI45SCRrxzkStCUmRRIKls5DCc1ovRhxj7b7
wViyEXZa2uSo2Dcg2Qgsylm6jgd+HdimS/adgLuLo73CLx2hWhRCPZEQv3tTipYMlKF67banGXBh
aFBBi/pHXGp5lfvtsyP9FIPCjLx7bq3TetBe93k9jjoNPWLDqL0ZadqpfPXZA1ebeAFwQW61R0Xw
WzUSq7IKgeur1Mq7oYMSwjqI2VRyPvwIUeA8jJz5TVBqfi3uWAfXgB/hR7oGLvW7iEMcNsdQS+/v
iYu5QTtlRllOOcl6y3qUP16O9A47aVUjAkOi1nIE0HBDMgJ+xXfsFRQSt5x7BhcjnXZAyAmwIg0B
5STJeLSUi3xNZ4IvmImAYnkBiTDQNV+8ToS6qFBiN67qWaWuKKKGon28S/0jBPezQgmyumvd6yG1
PKIm0VY7AT4dpm1MkX36MsQW3gSjvJwQXpcV0FKbgEnJsTMK/pYFXxXSqeMwTjk2zj+HMYjxQx/S
IRXpGgvA2A+RI8Q9q2djVo3bwvG6S6jn2BqFpXexiQyGYx0mG22zBdwFJ/n9TMRvN+HyMDBqS6SG
1YN9CsMQlMaJPa74SD6WUPxZYkFKLp5KZG0EG9eeXRbmbF62y386epyAuZrSWKyhdAGh2LSYe94N
WYBVXk+GjA7zn63o6J1uC2UziyNL85QonoIqZrdO8iwYpJMzgb2ZtT/iHnFEZuoDby5bQr5A6Jx+
daF8m14yqooJ3xow0U1yHnXOuq+Ngmr4Zm9uQc1SszTQQ0W2pvHD4mDEwBkHkIdTSXqI/AL18RtU
s702N8jhAsG8GlXzgpwqvNhL8pL0llQYZbU9i5EOR/n8nQNSjAMECVX5RGR7wm63JW0beSicpGDB
uCPXYSv9ow1PDlfMv/MqFYgj3eYduYSkyzmeWUQzJQaISyOFBjjlNfZKvK1+T6pBbhjWoo0ev2MN
0vN6vWnhKIED81QsMMQolwq9wd2byM5x4E4TZGT3pOuXu4B/l2jaap50zhPy1O1RyNZVkyVl7Q5A
lY6zULhYrQ0bYLmyB2HdXKxzJzJ0ZtAF4XA6MxtDTFLC05kEdY4xYjFLYhbVmiyHjyOK2UbEbOs8
J8qOs0vJbnh02uTPP7kWfAkSZIB0dPo+gvUX37hijPgRH7zevV+xz4X91zgOXGJwFNc4fSjIoUQR
ha+RDvmK5mv1Gf5AXRjnhJdwSempltNvlenMH/qjgNrKjDBgSe4WxRNzhBxvr0rEgAiA2gTCaYB/
nRSYoUEB7qGIoD0nmfFuuDjMWUBf9fQT4NTnelmXaNeS/kG+obMTQt8TdakzvFv06LDj6S9gWluu
HsXotBa8yHH5tGhn3N6ZawtqIAzzPiI0tyVNc775co/i7nYwvBv2ZXz5bHHJlllY/bZHdjXj3F9h
1Rg2HL5c8e+qAq3BZVPF4ySUpauVUb8h74I8T//Ow/I2nJBHiHlqPJy1TV0n5o6wdxoOYXV4H0Vo
OKsQBw2Xxxhoa96VmxoUBKl+RPyVPgal5WgyO8hDnq5Z3s/5Cm4kztQvUOKayhZtgkB5lHCKwXuA
elx/5uinLeL+AJaw7hutgcriD9ugnDDRLMpfIONo5dNoNZHa/LNV0WPf5nHlpq24XUEYE4hJADfP
Qk/PVatMce8TKfkvAib6mcmHTUH7LOhvgJpmjdilF5oaNB9z09l4F8Gtr282ERgjGk3nFTHE5qMK
jZ11xXeaYz7VSYgcPmJJ0WXUWz5N/j9jognqzrKZNQBLhRm6HLAGpQXWx/69hsKP9OCO1YNbeM3y
7LrqkaGfKr/z/imF78iFvUCIobr4BvhACkjT4EtDm5ZRTfs7ebwtyd8O5Gozz+jsLlcOAmh4oKch
W1X2Tpc5P7dD18FWE35HGxVeHS1bI51U0JGI//ULKjIrkI0Fr1ftF5br4l/7NdfTUEpIfFxsAuq9
RpgGAxBtzioLBqLGeOme0/K8+ou+6hITn9CQpgIdKRVTKvllgU+mNGeDwLuzsc5NRKaHLYlICHIN
Nq2IT/MNDvoEg8J1MyH0SXpcSJlkIFxWxKROsjmEjTv0sYv9MXbyI+HYR5AAYo3XgUIYuT0a66O7
celZSINueFIVWO1UB47bKKUY9mCKEI8yhBOAOw79fPKFGp6u/2UC55wBT/83klcM+V2ZxCaziXAZ
ECH6JaT3LXibLjG/DrUmwCJH+hImkdSx0M9/SK1C91Bx33+viXBTsQU83GTHZq8tKGmUf5BZY4tt
n323WiYiZTWC4CYUzkEp4KdeZsx1I+cPLtxEv2PimTq0LrcR60cIfgLxPS9GPY+2pt9DzG7axTYJ
kI8/Y1dlQiEryhw8h+cQ/sZM70FBSQKgXTvyePIzbEeh1i3LGptDUwe9TjfalU56mOrEUJL3T3f4
wbHfKi9mJsNirtY8UUc+0lNfhzTuYRc9UPY+ys/03W26KleKsurqyIdviwpn3yX9ZCuisiNLy2a+
/t9WehrChpYoCLwcMkmwuQFpEVAyfaBwWET1NeFVRGBKa7BNY3xUic9HXNqpZxPu157QOn/Yl0qn
/0yHrPhZnxNzX4owlEvLuIOIIMqntxMgS+zoaKH1Fe+Sj7YisZSRw1j8nw0mn7QXRWWkLavKVA6X
m7a2Ero6xR/5+HpeviOxddKAhoK7y6KGIhEr203VP8Ulb3NUl0YaIRZLpfLiKKmifewzuGEPhvBQ
HGDH+oonwmd9NbpAqKqQSZrl/MuLSDybO53ydJW7ZgGePAnsy0YJtA2FfTneyALBE6GmGMvV7rKY
9V1fZ4l2LVn/EhwVWADBj89rbhOmumEIWZMD/CofatKNG3oqX4m9RXHY2CX3oXMH7C3SyCRvBgBr
VRY5iuyIjc8nr0tX9thJJi3nCCsjAcK7pCrbOV9wOdSF8ZKGIdd6ciJ4gjMzBpGqKB+u+XGIAXuc
tXNbk9ywIuQsOb2W4pDkOWQZ+V5g1jOU0vIs3AHd7y/GFTRMnfYaWh5WQxYZRXmpIJhHV//W2adN
fbCuEvPGPyJJsSM/8f6nuVoeVW5cWryx8hsEWs4AnUh4x2INdrAKZ5MgxlfC6KEofS0ZvLV33MP8
TiEGUnUJlVAxkJo2RHcqZcJYKC4uuNnfgU5hVhBSd4Od1Iohwe4392CPhBbzXLit3zaDgI/8D4+L
IG1JiaYBgdu8dStU6/Rk1ghjTQZDq8cyDD5NPPTcL9Wdaf0aO+b9+jdnre2oaz+6N2QHfAh0Mcv1
mr6Xm71D6AdYeTrD11V6Jp3erTGQhBqSHhu+aEYe+jb7AfiNhdQ0DJvnoQ5k9eN5iw3Uh9UMehOI
PBjpVZkSwBn07d2RTHq7t8YFAMtAgcoSg4EKiuyVtzjVCdRuKpXnGCRYm2fhSikJrWDXc6nIh54B
z32YG1bXQu5FBBIlsD9d0djR3A5JdJpegAIUVOnUUKHqWZ+aTrCo4/Sr01NW7FqoFow0B+Bthdgs
WLxPicXmjChRPXOAp9KHEBe6rLhtrCiPsgifLDpSpU+g5p5uVJ4t1S0tGreSxurIuJaOcCbB/b8b
8vXG1+7vAnM8pJ/n8SBxbci22YtGiM/eXRVrU9l5yCVjqXSDEbVPKggwsnUvSbZGQt/ixJETChHs
3k93bzAoeVjWaZG4yv286uj6WDbuDhtR0ZIOBO3erPxUEDZrNrKeeuxZo+MMsoY3yaNXePcQntl4
vORjWHaabEYWeJdcrsAqLmxuz626Rpxudbrw1/N84jpuDNbxF6KOiYX2oy7pGoCy940NZs5cduzj
WoGPDLiE0BEslyzHOl6NQhW8v9pApWVryrzRU/ZMw4NbyZxM3fyZCx1N+IDIq+vH/qbJx7D4EMG9
sVnmoVtX1r5wRmrQpCFo9DHfcs5ZpFVx1P6uLmrOK76LMml3RQkr2k8/O1TzLrpM9/9oq/FiEbpn
cLJld68biaZgeJW35v8t0Em+TpYxzT7YlmjJKjTQU1l1tPS6E5ksKRqLiTjjxjpwGaOaSvnaZ3oO
+zoeWKBNMegf7+tH7SMZ4R8OR3porz3HI2txlnhaVtCbAbsW9ssxRMi64miorl3axTbpDILUYSBS
idXuMgpoktWjRSWXdv1nqaYqHh4mMdoPwoTQfY0UeEm+UxXuNxYYnVQ7REhmbmT3xoVzyMN0MXPJ
Upt1CP6JF2EKVjIOzce+bCQqpqlh4y0CGofpjK+5JQpzudy+I1PP3AcVSMRPHCXFYHGbpDVLIoOO
gdiEVYNCcA3RGwvPi7K5ym+7MlLz6DafCptKrZQ4pVAdXNBPqPw2ABLsn9kBfdgjJ41SVeHfsr4g
oNAk+reOsnXTlY6YD8CGGlCYO+Ovetqysr8lg+HJ0/ibDrgBFjGcGkDtQvl7J0gyuu2itDwfZQ9M
a/w7v2AWgsK1QrtX94KgvmtG3kjjTOu8NOnpyBgGqxfluNjcwirBBJs9HdqMKwpZ+LX9tUvD05hN
KG8f3qIYXMvleQxU2ZEIxeD89FcYFLAEOcMiWDe0094SprNWIlFPqn2iEOtfkWQqWKHVwj5Ik6Bv
iY1ZVdpWACZdWoJPW/M9MHWi0yGPYtQnRj+r+J2BxsqHjxHkLGcaq9atNdMfjnzEVYQX4DxCmNOJ
yALCijq+87LyR7BptuE9UW/qnOxjbyEprQd89c1G3C61SW/pwkhoJyCeLgedEtA1b5tObj+b41Uu
8eXVWv09ZTfqlPt+lXDhr7i1qTY+3ybPFWyALCtQOOGyYnnsPoU/7PLPrtSnQGp908Vrdk2n69Cp
fS3YfJoovxusxp31QN+XNO4kbxe3Ntktuucw+kO2xLD3TSivW4ryPaXD8su0h5tMYzgHdZO870Mx
bzsmfxGu9BWnjwAGt8p95P37wRXaizvs3YcKQIGzLvOS7XEPQn7DfSkbas62GXGwzCdCi9UIspa9
C9fToVbsAFPi2wLtzCxvhM+yiCq6ElFewmL8EGQiVQdsqJMMRpYwwGNiQTVx7CNziNfQGeti9104
59O/BLPhexOcMNggDSMIOIeZDaY5yoZcYxF5Am1o5+JjO7CdwBldB6de0v43fUpFpzVN7+KVMnX1
tmkOJEpO5GzTjftR8MKPXXusfviNYZpbsAbsybnfqH4YgKTckGCUnxij50wy3Av2cl6RqMywYtCm
ThLg4tlEyHe6khFvMP7InVAtTWHfejFOUS43grnR5QpZKUbwQ3N3EvkUwUC3zlUFV7afLRDeOA21
5kFXbb+Ox+jmL400q47hXqSQYcrjpUh1f+DdjGO9yrV2KHSjY0aCG7XQ8lEjmaWffqdsyKP8Ouh9
lN9nEtQ2gxWpp49BlO4DyEDPMre1/halBMLVpSOvBH0sU8w3nW80NcJHg+iUBTfte5sUgJHujENK
DF2gLlEAej4ZKtkfH/8XuTP583nwgcWq/8s2rtpXOqWAOI4J95o0104OiNNNrQMJ8ri18NIkF/LB
wHgKN3uz452vwmksJrF6/LBrbSCcVvYUcLUzbnH2cQRZWhbBR9DY8TGfDuCvGkmlmwvLkLv6xUJz
v9+3PIS+JNdJxCkvbuYUpKnjwkaoeXHTlFEX/62xCEy0p3slnQyiEkqpRiCwvumykj9AvI01k7rL
WtBEw5QPddTQHBZgNSj1TP/kT3ueiNvJfkrx4lB5EXYKVs28OkkTTJ8YXoJJN3whoxHrJtPXR8qV
9XmO/lnd5awyaqIQGOmOdchWfvc7DaICLWRoCkzLnRSV1lyWu41UTyFqWjI+iow+DPJU2WSXGLfX
9bsGOu5BeXkix2hqDxpUfwAKupipn+w8smTeFfPKw1XQ225Yuu/U2Li/4maMxI4u08K33uBrCz0a
jYbB9fIvj9iu7BwqVd4RMYg/15YANAYzCS6KoZG0NhcWNEqeh0fHuVehT9EYLNuIu9YNLNqIRJhy
HX2CnIHyZx/r801t00i5gBM4l6KhrTjWdoZUaP+bcw42a94lzL190IgW31Fm0k4o94NUKuRBhx7Q
pyMi5fn6RAcNi+X0e7USWrvdtLn7KPggHSWtgWo3uFRrHqwUL8IjaiXvMRxfeCowmh2JIe6vTK43
ckd5svvTj9OXJk7KbiD3dsE/I3baftuco3xVJ48ySVQI79lEWUK8TaL0EyUKpMphsorUht2OUYeu
Rxod3jPClk0iDUiB3aJ8euy3dp+rlzENOCNZgMKPl6Es9viEOYvb3VWKIvw2vrk1bsv3Cd/qLITp
R+F+bBWkkpp2ZhbjiqIoRj/D/uztfZd916Th0STJes78Xu1FKywk8tlAI1aJ6lro4/Fm+ZAp3ule
otZ4KtJ+ozYADQ3yIAwpHsJd8jJP19ZvhLkinyz8OM1qDvTHqtDDSq6MlDfCOZiY/KqcrmkwWgza
m2SmNKl+uXlk8NhixrqWzLpbAW5+QkGFa02yB+ZQQw6qENB0RpuKTWGzdNsUkRgTGllHt3ppb4PD
jZ81kVVQLyzkPsNZI9ftktvVa9GoRStZJX8YGbZgJZ/AC0i+dMVMhjR1HHkATW2N+hMqUC44Vdzi
PYxTdwjkyVHdw9fj0yPf4uSlhSCLVaL4bQulbiQuca8e1BXxbz5E6e7A96E7uuVBE1JwkfgkVbf9
aaqM1jahbeNOw5/mYX2qvFzqUEtN3lCD6pgjDxXfCR/el2yufOz8aZ9Eo4wk7DY9yoe3rCw5uRTC
Pe3SQpgtoaBloYmFsBo47b0bbHHgooOvp9ExWne/l4xNqFQzzv6+BZONm0HkPhqCJqMvVtn06KyB
1LSMboF3NDOs7ifY4X22GfAkXMMrNa05bgDClyN3dz0y5h13EAis9A3Re00dmw62izY/Ph51nfDa
Y0cXWtfRRiwb4CeT8LhwCufReZkDf12PXIgDKiORKvY/NYqQLQRLGSNdEupHaJZRKmH4W/PTQwi+
58y4YWa3834dIA2pONRE5OKFKAAoX9m1LgGxx2Oe4CFY3tCKNykctAHOrepe27euyGmbx6iGLiTr
urYoSE1kX5dFE8bIruqTMbdi0VcS6/2WfJcw2k8qHg8LWsQUVGB7B4Vfwe1FRCDu15jnpQa/TR5B
mRSBPJ1XOzfx9KXTsbaqJIGB0+9HyM/O4bGqLJL/+UQ+UAldxm2KC+V6N5iJ+lFeM9BH6n6WMexM
NbFYf95GKqtAWQu3egKmwCxmw7I/phSIGY8TqGwQAgpd6PIDnBq30yfi5z394IVnDNkI1qRZlxDB
yuARCVJ9iqUU2Dq1fYsdO5yMb38JC4QebjXRvPTl3a3VkDZe79xm/BC9wP1BmdfjevC3IFOi/hP5
Of7BxojID28a1TTEmQvfQ3lWZENZogzcPS6iHXLGHVN2MlpytHxFaBMNEblNpMyYf2YhcpDYlmoK
6/MXyNpDz1O78BcFiKllnx/7MdUXZ+CeJZxCkT0h9hE9olzphgiOdpIZKH8jNbre5iVfwWTD17m+
da62gkUm7N2U73Tr18uwILnfngjV6TjaZerCoUvtUAKpyEB7AfcMi25uiOU7USEWoykK/CD4BwcJ
4w5fVFGDn4Xfa5oXTRUSj3+Dm+fwMr3pc/XrdD6abx5PHWBxgoonlKfjcNRpgcVe8BnKfOd6hbmh
BLrb4kgwdv0P9c7WIbjA8ZT5fojAwZYN+BGH88l/erwtKWjiVZJSXWZ/LUHKrcub5KZhIOi8AYz+
YL8FrRvOt5SOa9Hl1AX5g9A6a1Uz1ynpkhkluCh4eyeH9jTiL2Q5pePa6DZyRIoGdpVtjrAyCSUh
+BTtPJD4wC6tgNhdHM+1v3IvwduG8mcOe63eolauaZGaU1AZoq5dgYQsgStZVvVcZ/z227KmwYXI
mRt9OiR+iQiWep+eSoqdEm8pzarLo6s61PEaijHGUlcFnqO19HEzxGTOlDFOHZW/hYS8E0hGVNop
V6HxHhK9z0m5Nr5WsPZ4fJY49z5naf11GfLaP+4z/UBiFAz8+jdQyQBrFI/m14rNK2dW5vmcPnjM
m1CRFy55/rYQAxtCTonA4hGH0wQsMDLmODXgB10Soe5QGAV0QSkD9KtvaTZOE0KTdMqjdAppv8TZ
dgSYSob3cNPTnM5CYqpWeD6U6f9X8Btemh93xVq8tWyLidQDqNZUtFZIngYl2hkiUcBkpWfqcKxh
RUmJj+XHFqnrXZM7R2+0GHykXb7jmKGOLzATcN263NdnM9Q0aYAic1xJs0U0HpnJrrIGu8OkJ5CM
+ZXWV9rdTPbm7MRYLpPIDAlEurinQ46hU2OBZM215z456CyB3BMiW8BTvPx8oPOBLwzoLswTVvrY
pkzqDm8CkxfhdLO2cy4wAneRmELAF0Kl6I0cpZJRl7jgTXJkSFtS6fA5wJ32kLWNVkBK/WJbot0+
t1tbcvGqIJe+KmgQrAE8yrQ4fhWjI4TK24H4hW1egpWRNjA9h1NcLsxCbDPtyhJbtaCKAF4rYLmQ
EtHxMBGs45HDevFe6AXqt8wh4FkVIrNP8EJPE/eeeoQolJRn1LWq3FYeRbFLXbTT14LPyG1/40JL
6U+7T9mGf5tj2ot/NY1qwBJhiRQ8UJaA0u/o5T9x2irSL4Z0P32joj0cFGQOu1iR1gKW9hxvnBQB
xIevYyN0gSxWthshM8U9/LtxOgfRDvmlrIKF0l3ZlTmc8PiGoeD30G8kN2QECspEAitp7QnUFjS2
cYyypYyqpVYrYNyi6075mGwXgMknmm3CBOWhNpt4xVaXkpdHpwrf1FTj2vuWhgIdfelb3JT2cZhF
mO5534sEvBM+4WKtVtds3qweJ7beNKnsWgWfPRGFHUbEAf4QGFvp7u+itL6ndThKHRGN/tvubUWl
ym7QDebSEGgtSg3e1FqhyJJm7zy31/cb8Ws1NM3PRfCrVApWOqa29gvdC/aIWUwcE2bio6+N4Ncq
bcTLI3eGAT5Ggb8ApPBcFDf62/dYDqP2avTeMOz+QLJyc+gqgVXq08oH+7zXf51wfz8rW2ezSjIZ
kAMffUnHZJm72qEARE0hoAW8Nf8c4LYWm/LgYtITGWyRz4z32QWNnByPGI1linPUOBN/WcF9AOO/
vOGiep2yzSlwStxgxTX1WsTqBdg0dznVcffwPg0Pjk6/BG1TfLRYqvC7PKwrrmIYUa8VcgWq7E78
Uzg15r/8AcPVt4j/OyST+zsuWQQeVJsTfyn2KkYQOyRMfCaqKYaI0w9q05qXxePSyZBmknNhikVU
ynD1O/SW4ysmExb7YrFswYbf2uesVAKwMRH6s/2JQP2svDhFdd8XcRP4wqzWazvJurSCLrluhDVd
jNdIfzeU2l/uvCjY3ZIrwINEvpfuYxMNFEeXEsqTZ2nAcYeEes9dnJtz8YsutKMqaaHDQA0efcBC
iXMmPzVEMOxwN4pgxKHGi3W71AblXWDICRvTKz2L2kV5kShDgLnTC4MJlkMuFZvASLCnNc/aCrGB
xU3jq9x+fcsHHmBzklt2rKySm0srAUPRzHTzKtPgMI96OmjAwAZlnJ/SCvM4EkycIWW5xbgRD8zZ
/xoK3I+9RKCaRW9Hb8qNw6J9EQ3nI8YkzuKaZNY53M9sYvfBHtFMQMEfwfKQykty05Zsi0cQ6idc
mJEEAUtvevyEscmAB4fqC0IwtKM2S6tXysABUl82r8+dItBikUqBA+NsDpFwaLFKMll1Q0S88jHh
nOZr/s6OfQ4yMqvYWCQf+qcBejs0OuK+suJW5gAsbHQeTqqJt7j/OQYKbscXvtvjdN0tWLQCuWbX
zMAwG23HTFOpFNdOie+SRf/gzee6Ntwrhu33oySqzNLzx4awzMrMQFv9QemvxYczP2VTdPrX1Shh
R2EGmyd5ifbhTDTVXYVPSO6FRJ0piWuOOoHA0Z3hk7JOMW3m02J9n53sasps+q0jpEbQErW4pADQ
9ByvlKDXPxCGrIdBBNfpji01PLPKd2wtFsBCKvUZ0oRFxoX4kqyBfmLzGSt3zqhccELuB5c1Z7ro
pxWVJMTY3xuS+OiDZcqUTPrzB68AYrzUEhMRP9SUoiYuTMx7I0i4q8fyuotjrA6m71nhNifK5m92
Z8zWvBOAiAHBQwNrXjCVInmPULracA4/L9erEeMk/dlKPSuNzFy8jP567HKOKVBr/oE9ibzmL5cE
fEyzXlzMa3NbUwJa3O1nm/KmkHS/jMigKUx8xvvylTDyMswkEriwtl68WWVGiuzVsYjibUSfWOxf
K4nvg3QgjV9NQUx+w2cxGM44mQaLulOrYShn5CTcWlkOTW7s/VyuhGhMqMVKvRlH3Z0jOQ6zE+Di
NrtLTnvlxJGLAD8JgvB1UPb9GVd/jwFA3fPsMhkF2bnz9uQ2IRvBmptuOElW33djcC657ACK+4KN
gpn4BKwJ5Mgnn3afUkbZlRsyZ3CoiVODUjFCo2jyA30Ya9fnnHbBFxS0XSl1k9tQhC2WnWm+2vb6
uK/7Z5qSaWFeG7qfjZbKYdDnocf43X+Xp/4yuf0rWKr8+s+p1l+/pwZ2xQiGH0ZZlrUFvSEi2Usp
cd3lnHhibW1/yGI/hzDe5QPI9hWL7PrCi8C3DeR6EyjDzvUJR3WU/Rsn8THPaspl2yhssyXgRCvK
fsh1AiFQdueLqQNmabWs6MScJ3L1z8bYfSiMpSbPehgW7kqRkRudfG2IiU24sskUi+ruVp3lPQ7g
BgOhCEzED31gihtZ13DAqY0UycTQc/iCv/64kFpAAHTIUumxjl62KdrAhHxkkH1TMbOYmN2SweWz
8epmPXN2f3J6pc/MXqBjC9KOt1iFeWcDXLYGTWHphrJktTdbFwQcP+iTZTIcc2VU2z56ga5Wzp4m
kuV4jfDaK852CYbg1ZgQmz2WurtDyYRruXbrFez6Gbf5AZB+l7FBu+2lMP0A/Ah7jaV4udFuVAqn
3tsMTwoSAS20eQMkEz7YwV83DW8y3koslp1vVpgK3S4ZdeJkiQOH9uuHJ61ki5b+Mm0MvYbWU05g
WrJ/VEH4GCHHkk717FI6L2MBbzbjeDpO7B5UGR4PyRNlCCDquwrU7zFye4lgbw04abjMpgMKrcr7
cCspElMz059naTzUPYAkZ9kDOOBn3krN8LZm3UtMdWI3v9Dd+D7gc3fs6XaCooe+pVvc9CkPVxWD
X0glBJyBVVpH/rlFDB035ESXojyK6fb9QRuZBzVc0SUadQO2Mv9+fpLKFr5Xf9TR5uh+15G2Zl4V
P2qMAjFHNiKGrYSR9jZPZhWg1CpFt58VDMC/THWnhQt5H9qtN8BqfyS+VkTwFWeCLr7XcOxtTX+b
u315w4VpQVwtKQ/xZhBQW7gk3XpF49t4jCXL7UJ+65pAwXePf4ODYGmNte+o5UmjffBB6HmXuLrE
qpvOeCZYjMWhGsQm1l1eH5s8DfasjO1Q6yPnCNo37AUWGOt2ik5HteBX1hvCR7EXj22PZhMZ2DHd
VacxiDTmhR9cTo3TOC5a5CKe07NIRL7JSp7idO/ZAdIVA/EpdU2vXP2KpT7dYRcFUPDzQYHq+Aj0
14bh8vXeD+R8EKcZx1KjaDRTGBAf3N+oe0bJWudrLIBjEoSfXwrEdl2qXgObUOUAJT3L+zbAccGd
Y6Y9ZKS3hvLOcAJy4Qn2Lgoifvv0DgEkbWeVLAJeiF5wPHvbYTdRPgLTxMfAS8UbZvFuMW3uwpTO
9l7vF3sNcCi11gLw4UrVzaukXMf9x3Qb9fLZZMdNret9/iG2IPUzru5Uq/ly4wbYWLPgdjcY5f0z
VlaEuvhnXGuIEuYcA9+PbBOqON5Qn1b0YI0KDPJ7F2VPC2wpnWobMbIVouTPslOm4JgzSwTl+aPZ
2088WwfxgWk7WRtzqDt0805k3v2io337ZWS470eFoSu+f+NiC0FSkZeutgrrWl168i4wwh9S7sDa
d3vqETffzo2EPBCM4DeZFQswtYM9xT0MNaKEb+3xdqLIP1SjsNty0BZROP9dIMfd9NeiPZxiVcF3
/8LvbXfhsEAfkESLFq6QnWQF/p1S6WxZgPnHIpM9CokHC7XucTLTiGCEOleRNihssSlSgqOTu7fu
qfc4W75QrMIO3fHUd79eAbTItUuZ2vY2FoMFyOLjLdMFvZCLzMIJBzWSE9ZQfCkMJ9nh6/f8exr8
f9WGAJt+GmwKMKQMD8akXhbEY2Sav6qzEM/RFc+UBj3xIJ5ZAUVNRUYyWQ2gGwRO1jvSLuK8xsDj
PYZda0y8Bx53Ir6lXcPI6bPG+NgQUWP1RysktkZsMR8ZrjRVI1GOzSMvy03swlC7YhFD4mL7GZTl
OsMt65v/JR4SPMfVHIYUoxnyTlB0ny68ZO4bKeDQJk71adDYLxSNxEdtzmhB+242WhzaqYPb4QpB
LtpOV84VZToxGEViJfIu9L3dn7G07CkPkn4i3XGjVN7l7zWwmaA6/S5w7W8Dr/2HsTbM7+GvR81F
e3S9HP02WN4ZsYartwLXPs/LG9HhSQyKdZNOlhdabuljJ1HZBjqQw0IvswuPeVNmfXHGE1AdHdDx
DNK1hjcoFGF1g7tiP14gdunpzGfSJJ/UHTh/EKMpi9vlua+G/K6GAf01wJamYrHlRlUQXLkWMZXu
AN0z2sB3yOOQpecSUpw6Fu1/Z6QtZFnIlKpPvux6YAKWC4CpCXDOWys52LDT0RYQiWqnEOF3fJyC
HCWkHBhwiG8zXqcaBS5Ix0K9ZXunZwYbT3SGF0Ze4y7GxPeMRCCZuf52reEbd1EQuAVNg1r+RmqZ
UNu/mnxQVzS5nZONbvjzNwyFeQUa5ihtEleNq53YjUn/wYzAmwFiaulCyLHQqGZQxE55P6evYDwh
gUwVRKnnz51G7f0ARfxWY6TnMtiyfU8GUJ8VL13h0Xmw+A0Ml4l7gprc60CIY0Bdo7uVBL0NwHt9
T60yT4E4ohyamlMy5JWRdtmfqDJccI8E5uLeZ/pmXpJnnRw4Ik8o+4o1E2kDcMHI0BOUuGY/Bfh2
Fzfr//VVDYIrflAXG8IBw+vSSXPfsX/6AJGZdE660C2leiNawIOeLmGLbfmOksX4QWA2JN6ySY/r
S3E8AEunoywINmzTAFjPIVnu+OtH916njLUOmqDiJSj/ebkzeTd5qegOkSwbNr5NTjOVgynT7bkD
NmoSaptEfUqzbB3RdBbIFtRb7gWuWAOuid5I8nI1FeaH2rkeCdDFv0EyFaPtO4UFXqQn7DFa7Uin
p1RbEaMtW99OCiAm3z/5vRULnMuFNgWJVSvYBZSt+MGPOyLCllRCINQFllB5x1pGfVc7p34QrP9C
fXFfkb7eOUL6PGiLSuBuVJG0bBeXE5K7ODTCdX37+MmTLqBVPW7h9ZOmT9KenmbseXfQNmBeBZ5y
+SrHopbzNLtfO6tzv5SuvTmDfwsD+UId7O1M+2EM1Cy1oiU/fkyLG9DtRF8t7IGCspszPy3MpDcn
uYl8UF8LFB94f8gw3/XbEThiigV/m7RSZLZSRwKyHyCrC7Z70BXIwsC8V2zEFFiuMDD1ixKM4njv
kiOQsgBFcvA0sA6cg5rE4UHznP8WssL6i0x//CQd/uJOXujvCEImbmC7bgbv0xM1N/O+O7t0nBg1
KwdhtkQFAfOX+9jE/9JZavIpjFQSQP1PCBs2sApRWl7alX69UqnWh3Vv+yrpFa2iZ88mYseFqB87
8stPWOGA1genVgRKtqEf/ks99m60+cZ2KWKQ9uKCKma9HqmgkZodE+PWJuCfucfWNzrV67F/MuT3
LQp9dVgrt8zKINqmKanj8KIrMET66i0dv6FdqquMEc11wkDWrFbHDeuuZn9DpefmBytlP5zSO46a
l2P2TYrwOHtuKhLA8b4o6ZFszFD9jf8GRq5nZw5qg2mG8k9YxDVg5nowkN8TOZnyxv3XPuStZqCw
xklEtRkPXWpurqw/OeSCLWZcNFEMYxuIDq7MGnGejXjgs2zv56ZwS0uxB0chchmH+V0E1TgKeGBg
MtNA76bp7ZM4LTEaalX3Chvpp8rD7vrS1xpa0bAdgmTXjzhWBo8sb20hu+zxfwXAeahbVHIat5vS
N3ThQwr9eGtXKLPjZG5R97AO6pWi9CT09qOrSpGS3rJIzwCaSUB+hC8JB4siCxWcgbbtndb56QAT
IbLXZvuu0LjuOF8QssNhJk96L2EtSz+M9Gg2KPJMM3OWiGUNDVHbVGi1PohLyU/0/E28E2D+8tyN
farBbrN4aRRAERrjZghxUrt6ekMYeoR8G+ykaxsKdPGKe5G2Q7vf3ViI67sr3glmwzvSlnnumZ+D
CsdqsXSdqFUxltHcOrON5fHoDwCJHUQT4Spc7auzMf8HZOXzRm5kJfp7PE3nB/SmP6a1hpzrWlZO
7HeLjSJQ7CJ1IaSunnKZAaT96Z0UcVp+xLdkCpZ67eKhCv/5ZCwzYorkGLeBNhHGYdfhyj2WRl9+
bGDNLSMF/mxgPxg1NRT63qNcPTE+9RdQLaxRSW7vzvi4FYh5oTGR7cMVTpEuCRHopO7WWiXXuQYR
rAFlKfdcpOndgEY1ePrllAWCyybrqn1h3j+9bz8s7qkRtgFj3i+sFIDeJK1KxOPv9WfkZMyyqQOP
UnEG5fHmq3O7v+qCv2FjxCwPfSlqnJohcDemH5E+gapt2OzdYmoKYxnGCnDCq6AhtXxEUbVM1ODM
JVARzULqvVqXfC9NrN0YtUvdAn+jo66Kxqo/HJdj1ulds9Go/YFdr1C23N4uYHVgpLJTFbXs5WPe
X0skjDfHrvzgnKN4Tj5IYmbe9CEPovzIQZOh+PNrjOkkeOlL0cIhY37knjI5hSKbjhZmF7W0nW1r
0vcEtGvElya+qjGgHdyy0TiqDDBJNEwp7VNvg6B4hrFNrbDIhS6peOMUpv4ZfDX/+E+Ce3cQFGXP
VJJa5j4LWKybW5x7Zn6gvJnJekCMJu7aVrEJ4dCr/adrWA9mZvSdSAmkL5weK31ZTSW6HgdpVd1A
fgg7L7MZfACq3c+wxXItHfL5OcetUcWzs7udJ2D7dAmYGUCzac66v06snm2b5COqG40iGalcINVB
g+3V/WJP6BiC9GTHXeHDMN9K65UQ/mWURlGC3Zf3Dj+o3+xIwhMh3UtiSQy+9g7YhjHWw5JkJwwr
gSGy72VkwMR48l0n7oGyNLnNyy9FRxGnD1mggZbX9ZocUL69NzygYB6EXRz44Xu35mp8UQNU/YKv
d5gpSVVifp+s/zIMHkNHnNDi3OX5hGpYdEvKb44Yta+mDjsHsZlgt2bUeM9I1Ffi2MhOJqdckiGj
R4cVwnnHaZCyaVcrshGyHDua8LnoOz57+nJD/1RpeCstkDSAEUnp8q9R1q4Ob+7RSoRkePfwpYaA
v0/iYfPtKEIGJydNtBHLIxUIsk1PDg8tnMpPxaKKvvyMiNAzcI/2VXlds88LQYAffZ1BWOOa+tFG
D1g5Q7eIkzEm95R/kPErbCJowhsEKsfVabrKcsEtlo7abTEtNz2VdVJwxJjHbXvauOxRGqPQRAOR
eM5P+oUpUwTAQNWksB1RjLErQcnoNgZRIJJoe/mtPy3QpsTm5sJFc6ECTah5K9TloQOVBbsu4n2G
gFc4aanmDYu39LpO5dYlZpmjodUno3U8j9/1pPHP3PL/ojpSLdfw42AALA37p29kvh3pj4Do2Q0G
Kz8BknUitL3gvNcQ/wxGp9i15wyU/At0H6XGvJ+K/BdjvknTGa1pbmq8M59LTZQ0XthbsQTH2JsG
iZsKCRlq6gzxkkfar4/saQCv9rIcKJGkxiDvBifq9cM41WDcP0lNliiwfObgoPTThfZonZRw4oQR
Z2ojipJybQ40/e3KcLstVXqSKWWrb7z7Fsp53gveL2m5I/rSgZzmQec1dTlRU8SPyzSifNuvCPoH
GYzw7/ntpQRZDmI90HmVsdVEn3lF2425QoYoHRDW+mSrMdUdG/ojPT0uROnDMIbFYohWyz5ChUf1
V/icxlduCfgxWj8B3dQYveHFjgOgbSGzBmhrdL56zbx3pGgW8VhsUPbKdYGdnOv4mxnGhK/HzWkU
fbQZXQfmpcX6h+8B+nMv9/tSN8lf91LcV7AiL8c8SC6/cg1Uxk5j9LT6IMFlnmMwgT3+P+udYgcN
bUK6gtKQelCnvfHaM2gzMgXQV8m/5CRmGxozlFp2JYV5HLNSAFysMxTGvZru9QAqlgr/JGaq6qn1
AgRkY5bdWD258HSsJLS4N+kGesWFQNg3sukZQd0OX01Kg0V2MWMd5tMggAnkco/YxI5GezJaOSE7
wzxZzeGqaDpSE0sQkrVbOXOh3nBaxgbnWpvzhngALpoleE1yYqRJy5XyHSldnhYx0syZvmrP6msP
anyqTjAJveWYw+Qipgj3f5qXAmpqRD+JOKrgfuadR7YstoIxoby65+ooL/mOHN6eDVFdp6uPJvTV
Ei78ZMVc+5QToecrqXk6vS43VkQ+glmPwaBokQtpBjK+GTBf+r9U7y/Rui4321/JucvUxBKV/D8X
Bj4QwH1/uZydBLWpgeq9FviLgW5lBOW9BUcWub+aHp/0tSPnYBSvsfNi53tF7sDrxgy7446gcUL+
49H4Z0TetNukJyLb5s2sWblU8VKy5LxlQFjmrmOLyCbVV+Sg7gHutV74gXmOX3zGOKkQA5r7OG5p
fH7a3j3zyGGQsfOb31sAFU7sQAlJF61shQ/JSBRVc5TZg5Nc3aWdsc3hX4o9Sp7gAdBU63em06w+
Hn0W+RNUbdq07aQZ84xEs0DDUf+6OvI3SMF+I2EJ5XLuGAoTBqqHZn0+1xYrdEOBabgI7zd5ddA7
s8MH2g3N7C4y0f4Po83nCx+l5YXuXiT8V8XjR+0kwC8p38za2kXEzuM0BYHQDSAvebrKPyvQ29+N
J3tCQJqH/GPMUAlDgdcUAdIz/e+f0ek3aKCgFcbCO2FOsG1lftdlokN/tAYsDePUeC/RIK83Grtx
ujNL4PKAZyrkgFTE7xyJwZ8UAe6zXUj/Z6mdgCA3WNInbaONsiPbVEU8MjS7sqHqbHuf53xl1Cow
vOGF94ofUQQNe759uWagIUvQFIkr+vGUDs12GwXJeH3bEkUy+DTm4F62COnA0gBNgvgNwcgE1cXA
3fceV5k0chePinrEx3MGy0sYpUsKDpkzXhG/xBfLfoGU4ZCZoHV9aAGXGsnV6pVZRoGPGXMGWR7h
3nP5u7grQr9Acm+Kzj1YZNo9oLn1jS+633DoSg36GyvIGdDLFB+TPsC+kytdkXfv42ILkgJZPQEz
0jTUwbw0r3iKA7JiCbktSSDQVYIjHr6GNz0jWf8diOuznIHU1CoebSEzj51gRKkAWkL6inSLKnsI
OlU20jECXoM+X/NqEZifXsAe8kT6saSRIHftJurL/mAYuJfrDpDLe5esOEL92w1V/GYH5sclq6uJ
4MA5L/dX1usQmfD3R4/uuhoIVcGzGxGzH5++CWB043wzH0xQSCa+iDAdVpsLufk009xRrfuIyxyY
AO2fvTzT3La4cWzHpgvsSmURTgb4RAYrmUN8Zgks4qA+j+RTCCQzCB/PK8RvJAJ/z/ytwk1HMe6A
H880yu+FvL3OI08VEtfYTM/ueeXYpLHJ+r4xPGqFXpgQdxHU+moqfgbCAfNtmXwQnB9weq0o/OAH
mMCA4nqXDbhlDuIqgVAidVPj7XxWSmJiTKPSXtm8gHRsUZSA3Q7l7iKhq6HWr3qYWcSGAfjXPFct
4xb4yLhLB5YGqFqlfLMygHwL7kmaUZoeLdaM+iGj81JPWOMSl7GVHKQpimdfF8NL2IGJ7pu+5l3j
UIyHOQNNBm5mdfhdLZX4abmvHu0JFb83VmEJu0kHlx40F/FOcgfzspbjay9+nVTgRSYBC8DrfMc8
O+sFdT1vFkv4T+OgdF4ZJkNNb0OmwP8bX9ljTBl057x0Pqpqbs/gWw9IG+FKugLyAGlodttGdkZe
dUqEqY+vaXREFZ5A4GsmO+WD4gdoHkAU3zV4aG5SYb6lTbTDPQhE+DopH7wYf4VmsWToDlVHSbiD
qdf4mQY/qneR+ib1HWqKjaRDiKNVqsDdO3wL44j6iCTTQnYS8UqkEOU+IaU6QyDWwqdZBFViBOCn
DgYDGO64CF+FK9fwuYoiCZGGZK9fBg63+fUwGQli7EAQEVjVRhyyAuZXNJv7lKesZZrNb5gyYANx
7i5E4PAUZd5PmDhr6oQ7aX/so9LX+57B1b2fQQQqNCnEaF5QZcyvZ/agW9uq/jwVene5Lh+Sri1P
sLPVZHwPWoe05ZnSztmEIR+3VV4aIf77YNXPaYBJqD/hjbYomel7Oc1jwqQxAn04yrEu3lmL7Rt3
FcmSYa2PEQXZmuCv91b4N/pql0FAOlgRqhJifhC9p0X3bBhXWczaiPdoQEtPvUYlmH6waHDA66JH
S19tnCEzc7hGFcxOtK/JfEOIyL/SnYAkgHDTvz2Yw+QoE1X2H0CmNJfacRLK8dulWaCQjXfspCRV
SOwnQRWU4lgdFAz1e91WjNJcvQBZTK18j6rEpxSSo7XG/wPFxmCArRjPpA2Qiy5ZxlPikT56yMDg
OrVIEe4Y1FfgEBDGg85nDcT/GqYKflgdfYthEWAPFDmlGJqjaIY8Ol7wyJBM5eEqVtpleqWljwED
d3q+0/Nbmqve6Rib82mGfyEf5eslZ1/DgNpNne/+hGAHgmnllgfhgZlnUtsHgFxKz+FDto9zUSei
DtA/Nk+fgHa+eBj4y3WG5RfV8sQpJv1zgeF79XnPKSfzo4+I6wdKb9ztsrEQuJP32BQ/ptaOBQ0h
gf+GDDO86MsDDsAmjfeYY57tETNUJKtiND+uGmcmT2l6YgkGvhnF13jJwT4jEPB35KuOmajviKEF
jzUVdhC+muFbQCBUBrX41x7wzj9t9yUDN4DWTZqWXz4sdQA/EwlTqJGCcZbVklmEELPC/IYgiSdH
hAMAdOb0aS7xd1rf4VhjV/xh8xayV/yJc8nManzFFAF/316dRMK587lwU8pC1R74SdsBmRSHRy3S
nUXMSc/itE8RUxyyRQXzx4W6FxXcFt3cGyElr4KN/t6q+y7WWZSc7CXYYVTLrgLuebTugVgSrFdq
HVob2I7wQ2thxkaCfJLBKecbeDP5aOZoW+AW671SSy1CRSTfw9jeLrquY35I/MNI2I+nNzf1aZVx
FzYMcIrvwYo4KuqUtKimg9pclG+Vm8sgO54/KExZCV+fXTITPUtTxay4BSfDqVEoOMSDgLuEvndH
+5crcEY7wsBDKm2iC130V9TphCgonDDf8rkIK54hPGeHJk84jBryzsIgepOFniajPZEa8aJFWH7w
xiOMgg9whuo0QZ5r/201MFqdw1VLif7/+Q2NkDKX64WDZudJrLr+0bYI9cOUhG0IFqr2UfPPJZ0t
C6rs4QFgcQFFTL+DoYldLFdSu9ThkiL2syNqeXpgJn38k26mN+p6AXDuxjhc4H0IcbIgCNhQRe3c
E6j0shkLLiyjs4STyhtCbsgldw5HZIzc9CFOqC7HAYxQXDcBtjqQCtheqPNlVUkuT5zQ8ZwSnSA8
EBI8RfFkuch3FGskd4flJjmm2uxbAad8WI2OylSb7VG9oKEdHSCqDMMR2JhHMMnNBUrwvroM1mQ8
CRelOHb/yeq9feOsbur6ULcfmuY5IRphkfUWFG8ukOCj7oDt2IFRBFoRyT6W1LvjxcQMIDV/7tZa
5eMQHJJwRfcluT9sbyFZKReuTjCHSqyVbMtvibgSLJqVf0ONNtsgcr/H4+OGBO5mBCIGMKJ5aFKA
OcEs5JYrdpV0KGQ3v1X1K/3RrN09OgXs05dnJEaWrYd2PnYvZc1DVm4QpzeTT7SENHNku1F5wcYD
FAUbjjdzzUAcLBxEOuffZ2uvF7ra2JncUb4X6oi2kgJXlZfflxY4UtIc5cNSrc0DyCT7XGJkdby2
pO6CyqRofNNwMghK3gA451JYxNoEfYPtS7UQV3y/GRBNCY+GxUbly9TP74mxkWmJLWWhVbPBlAfn
chtESVCMZ2njahMRArE95KBihWq9dPX0L4XMtvS5NmxrkcinegcnXVk1VhCRNs8pXFvm28am2ycj
oyeClrJKVB67cM1tmFtYrlTZjvI8W9yAFlOwOzsGe42c1ei6sFWuyshZyfS/Xdc7m+idFLR92omT
wBId3SVGlywDzcRF4Q6NmPlybTjKvMzsqLugdCFNQU7C9dK/U9IvFSxDQ3W3/4lX3F2ROJ4bfWEw
tFJXMkuMu8A14rC1XfT0zMBaHGl0pCA52P0ACHJ0qiOW3lrT4ZYSk4Svuh6j9fnITVcFWa2OVUno
8TRNbkDhz09fXHDUDvKDEb0AGxSK8ImUneYjMpgyL2NQtXk0ejlXYyfnWptPInRPLBnzeuV7tn0x
SlFOq6zL7SyCAPcDYkMfXBX8zPdGxUPM9T94H+WE97lZgLclhLl7ZfQukuqjwY1g7dhVSJ9A9jyH
2ahBHN8YY2lQbadlFjW09rxo1ciJmC9L3+SnNLHocYVIFctLmnc2EICUjHZWlqOcqSvw3RvrSuSB
SmzPN4l1qAIGnDIlGKA61NR8T2kFCZuHdLKOfJESwbazP26Pwo7FdQTAWnU83zjok9KApkcjnwOX
dweiKsSL4TbBlxHHuJSYei9h57g1sBuZaj1JQ8OLLWSbmFbIGPIipZ5955UV1u6KRWVRlaGjWl8j
aaIUdsbvmUhWClcv6bkJVGxoXlIP3IdTqOHdH5lLiQMxMX9XpqZDHtLgINbmxesRxpjZxvf/+YnW
Z1UMSNaY3sumz8VOaAXD6OOND+OSOHiTkkrQns30CDN37rxcqN2/UJ0d6v0/3CHywiaDNf3phXsH
sKLaW0LLR+kyOiDit3Nj1PDiofKD2ZWEGXkWNpiyq41vnEuKrtRarNqhpMa16prcqJEUCftce2mv
mvxWtNSByhygsWvgUpqXgQPT927X3Z0E0lAMMEm68eqosy6g57O9pmOtsisUyCo9WCUfzeHJ97gH
2DtgVisEXqq1C32At6ktQ0DhnrozX3kDJ9wBcTzDpB8U3YBs9wAwH2JKqcr1JyXyMHuVqDCBHd2a
4x11evcpYz05J2lzmt8UOdgRw2Sq8VIdiQAVQ5Mub4nUeHhYEkV3R/TB3yrkOdFTfKNShksP8XOL
DsRV1JhAwe1OPMxOdTRohJqZb2zX5slDVopDpkVAwP6M3TYGis4uj0xn31tGjDyOEejOreUArTKK
EboJaJfmPNx6zEv1NlIU8Ffohcmcv81kgc2ZkgzZ9bH5WciIJ7cLOHeWCqItub8OmTLSXFOUmh/q
Qv9k/kzvNZACnYac8BnwQvyEqVcD95VGhbwa0bbf3FbxzaM7iS0hpdE/SqHG+hnA98Ahvbqvgh7X
U5Dj5BuwITpWK1fiX1gIA8oV17/WbGMyZZZ7ChYqudeWJoIKpi+ZV9Xyam+E9EtJzrrbk+9AKIuK
5Do0HOkxyF4j7eJEAba2QwlK6x7fl+HIJf1iGf2IKJUqonxBWR9nIOaCgHD55V519/wNK3u2v8RN
o788fzIj/xt1szgUMR96gaiIcEvetEkaO6E8qTLertLnpGwehbTHmkMbzd9XWLsOSXA0LXG2kZu2
XPUhtPaSxIi/4DkmxrwmlHPiKPkH4B3LY7XEuwlBMOds0hfVplyf8ZN+Ix1Su6iRR5K4XHeT1185
UFMarNnPzPMlXYyvv1ZHjeCiRO1syu2sgrHkwyTLtEOOE6gFToQettJoVgzAILoD8x6fVTylyRw/
aXPz50nHAOMC/mb27O3KcHU7In8ztiE0ctmGu7OKT2gj/fVbk4tRulCVEtw/KKJh1ygK+3BRDpgd
Y5HoCEq0IG3s395zNAZjGO7QQUiBuXZe31G9VMrjk7aY3e4DEe7AkLjvRdXc838ah56Y3W8VSdk0
1BbWbELLK7Ak6LvwIGSUZcGkHeOi5FlGxzNMf0td+l1oqdtpGGwnApcC+tst2deIIjC1B62L2aDL
wHYnU1l+jgxKal/oLNBX87LZxnU9+5ZMCPFIaWfPqSxBfHPnOWWkxEeDEdnNJ4lJG77jWLwgNRvD
r/69r8OEA/ZqANXaHjPDCXobW9L10T05aGOptUrLy1mrScWJH5VFDDy1yFM0QYE5VuLEOdNJoeRc
1WY0dO10IEvWCn+5JtTWeoPHSzPl7+Z2R09VbEhSqDOrr7h+s3TzBRO++4jYGn1rRbeK/IHRmZm8
k2F0oS+uoPdPEvZFW1tefPQFltVraOp6Gkwy4AKl5z3NWP4tEWJ2yqC5F5QqlxuW4jZxsITtOHza
Adw6YBulUWSPyG4pNGgBoz/Fl/MDNpxs+C6qsEQcniMv08fH+E0oAsoIoi27LmicPGNBg/6uREb+
nbXgYwQf66a2KT8+qBWt7j01G0jwQ4B8cktE1aHukAM5Pzh/pCAi0g8/EQ2PEfaWokwjHCh5y+jR
jgGG8mcMyA8uOPOrdKEeL128uFvvwAuGSN3oy2GxTE4zZmiBDuf1mEHPHCtV9U/KOTZKWKoS1FKl
cn+M+FiEMEAA6HMegfgxyM2qASOy87m8mArcA/zHhWZe+vRjx3GHHRg6hLAt2td6jCla6KGMqRtH
mRDkqp2VCx1BLf4Cyde0qWbRlj1Km7ykwHnRndL1lN75KEVIELpMeluuCado5d8t9wGn102ae0OP
rSPxZ7DIqNE0Zj5OhswmRKvaJsv91Gck85jzKVeMBMWT26GfFnGzKMUHNV2eBhKtqDbNGqsYhi32
NnRGP08aTWDjEiL+AQNuXjSit4x61xZ8pCgjz6WPmYhLWPHYrRobh31DfmLwPHYKgxM39f8fxvN2
hizsRzyDeB2z0zTmN6SOh3Qa4HBLPL27jD1NiLtS0XREXWtGba3KC+9Lww9ZUAjpjIN9FU59NL29
GqQ2GHpCdNvlkxBpc64mGgPPdmJvNuFDywEmE0/nIuyuV3b10uKKLWen6l8Cb1xifGlydgHOPsjr
qfEhFZ9al7NjGSsJcJ36c60XqJ9qFCH+RqpFy/TlE4zKpZcCyKcaZAc6TaP+g524LZ07ngDSEa1y
ruv+Bsd6UgLhg8PYZSMSqLNM4IV1GubOGtHvu1dqAPgA3DQFIHKJW3f0SS3UtYJOFjyHpc9TNHBH
VAGTnvo5sIlvB3lS7+3Y8VT58H++DybU36gAOKoSWqOeL0K2Q/nmh0KSNTOHfxNPTiJ5+eVzPrrv
uFgE8X+izN5axsaCJ5KsYlm3VDDmUZY4fkFHN2LgJA4fBpcptERZTvcWqLKU9YqD8tEJmx7/3OsS
AWozKt7/KPZqP9mffWqKYNIyriqb/BBKH8SINbw4+jWmEKhv/WXk53b4zPd+kWKzXQNesK1m3lFw
gcTH36nT7uskSC/z1qBvnC3aCF6vt3fuhV85S3T428i4V3IFpXnM6jJEYBnxiJP7fO/jp1H+CvzP
PnicOq++/+jmPdTQ8/5rNB/BAo8rWAR4v7uVT7ADKXnTXeF8XzwdMehZ9a244PY+G2s4cAby9srp
UDTzrUfcBRNxtkOCLE3n63/XoSL1MtAFHh3ZtZ1dPYJS75m0nA2olOwEWN4uc1IMa0jBb0skZtcq
z+kGjDe9t/AyDybO7moVnTT9v5iAbfMYvrLGEe4Sp7U/++DyG827W9TMn1Wlg27ITB3zhcS09GTf
v52vIhPoRw0HZHj3TyGT8tmiA3uWYJPeNt80zE9i7I97mmgqIPZSOyV4edM1ePUfvvrwe+fOa1IZ
3i/DpwMNhlyI1PzFeDJTxdoe1XjKkNlFqied+EhI8vOg63+bAiUoTTTvNf63J9SWL9HrZhbuphSH
r2mjfNmA4jIJQNoOuYqUxgE0F/6DMQGsOiVfvM89QV/rtJpFgml95rlkfpy1+Rl2Gl4io5k25XKa
QOVeSxWKp0C/odyUcGFdw6yHSMBQofUgUZyDCL6Bnyap815d22R3C7tqlpVwwKmZPCLKSUSjVQu+
2yI14276UaA+yTKQfzr2DuSl17uQvJa1J76pBivppnY4tgNUTP2Reks4+FvbhiZ4jwwKnSwoutFC
mEPS74Ntv0c3IFLJajiT0nlOVMVyyRx6INnNTelJXJCHwRjbXbKp1jTOm+UN8dP6M3zCeUjDiojx
f8Ned2zQ0RJu2khIaXkJRxQfNWVHzWcKwYLmF5LbmUSYGa2g3kz5qAFAtup7npPKlMpVMh74vaLl
4ofvs9EebPdQ710mDIBpcta/nWHYYpQ83Np8gy7f2pXpVjtFWzkG/5qcOjh4V8CTXD3yvdpwzlCn
ZulPNVi+a0EHXLa1s4PdbdA4CLcujbhNLeWyGTewU8RGyDfsAFbSfR8VbqksPvFyJ/fp6AdiIiw+
Ux0zSE/jwJcndIc43K6E+CFT/UrZ3nU2tT+tsw4N8EZ1U+9ZrX8RxYeRp9tErSLxKMJUU2UmSxwh
wCJATKNG6EFVtcPEJZ9vVQGg/x4TMeMf+6vKOY6V45PfM/hLNNZfNS3VY59e79ZzVnOuZXMjOMkn
yXS/tLI8Df4e/lYI+Rgfp6HOGE25mnLsDwk83tHgn93/mTyMtHZ9Hgo4qbP/I90TeFDsljeOSuLE
Anwa28VAUaJXjx245IrNQksQakxG1+YxTvc+CwqBOXVVDgAcyxPE3Ky+tmJIf484ZQjWV2IdboUw
HNWKQpqgJd5VBR9OSZKy6eQzjbg9elMKZwxxXOA4MfKl6vF2ZHRQofh3AVDMOBi6vSRLiuEh00Vg
RuvObNrrED0xiWZEu4oRyB+F2LEZcXdfuZ/rpWIzcHuX7Z7tmCFrcXnJcJGHDds3KgxcktgZcUD0
unfamnObCMhMFBoFc7nqGlUdSU0jSSvizeGaIoWeyb4mU2EikyicP14xuwHh/fRp7D0yIc7PZpHB
QVUXaDvvprWeBRWProM/1FsrNi9OShjx+t01rTQ4uUfVLFklrhApWDN8vM2C3/G5D/TXu4WluYli
7LbJxvXkXTtyiQk5RQWfLRgEfTDbAFqoZR5EhRlsAEXVx4Il4uizsRJWlnG15aku5li2atSf4pwl
dOBYRgjACffrbmGjybVhbg7SZl3J1KqnCUFa7jMOv/aSMIJDYFwzEkKP3twO+L3QYSnnXmPpvj/C
Uaz+jWasO+9FabK88nhoGJ+esZKXTOa8l1+x+Sxlktm0tLk4U5M5U2oHborY73xTyTsujlaBpsQ0
gkk41GkT47m5JADhsWi8wa0vbRydkFTJbq7GLakYQF0nvonvQ6+2ETlu88nMtlpdQrlIOYsiMoWC
BvtC/oEf3kwBWiwAiXePqtQwfTnLW+ZknXdQATcUkbOkwC0qXCdnzMHPq0exbbSHkuTmlTjB05+F
Dc4mvAd4PnYuLD0zcHVuq9ffJOZvTvGy1djo62qId/nZ+BDzuvOnzQYRgIMEjJoTRPw06mMfmzcu
M0UjKE6Ar2s6/pQvTxs8bKgmHtPzdKCe6KskWTrI/qnULI7OLEwsaItoDFFldQL4Nojx0nV2+Pav
2do1aPcqdAKgq+8gYjLpBQ0jaByz24vVTVPVi14VM+W0qAUyPpR9KhTRb1PrldN0CnKP4RWWCJDY
NZP86YecVWiAdIfbpSPIKX3AZcnuyR1pS25v8SmRZm7iH2AuTOgX2ftu5z0ST8Tdb/fsgYlv2cle
3jdTTXrHFzcuI0zJvnOnPcXxMg8DG/d1kWqFvA9psbshO9e4dKfhU1F7xBIRMTkwwoLoaVFPPfB9
GgoMDilZyQTlhVW3zKelLsSNmfYVi5jdB2GqRVX3KmKDVLaoyhdOwkiXNt+AJcDOFWLfUF5rxWxw
zturjjIxfYJ920y+Ldbb3QyKcaP0AWyD6LhTs9P8aAqz+R0meqCfcwp8OWC1VOn18+5XFFnTsZch
awBNZbN6emGdJXxqMYIteApWg2RMernKUINNjzYUqthmIWspAbWdsAGgtqjJyDUzLGsPvJIDL4ud
TBfG3AxbWXjirSgfdB67686JfuotvtE3GMIitb149PlyE2hwj0dfvXZh+e7b1C+Ae1eHKYfKi1to
C2PhNRdZ62cfuFf0ElgA/LTh9oa0TskhB+giHK6JomnTtumBBpNqxYpFaOOODHl/7GMrtVUjD3U8
UKpWhwIlVZjsIE+5JVxIOUmdirew8ckrLmC3ztsvuUImPCli+hx6CKCzT6ZcHNqTzGRTi7fHvsfD
GouDv9zD+/+djj2/e6Xw5B3LhDQSWa8dfpuSMFo2y5EZSGIecSWQqibw0W5GVnoMDMWifMlIJxev
3X8Al+G6/gKgI0W0JzL42IXHmRNlytEQ8F9gI5ygbLL5UCkSHlNPjZDEvkNwc6NwQ39Oqo6Sjau2
fLEK+O0GgHlANY4TF3voqD0z5d0y8ZVTlHi/wN+DuS1TNXM67YOMiKOjfYhks4rNJQMpKZhVG8yQ
NC2re13x7p5cK/wRjjcmF9DkjSB5O0k7omyYLLtyl1Kh/hnXptQhRbNdiArwmi928NpzGv6CmGjn
PV78m+eQIpnRxNcbwoQVCFdfyQhWXfOFk0PcnmYjHm3l7JbURzBoNnFshX7Ro8a3U5K2zn0H1GTD
Q+ligjRASRvCE0Kx+NY6k9F6/gLmWYfG7zzQn/9KocCC1SZm8yyrAbg7imm7SYBYdTOYQmYLqLOs
Azw/nNl/9CJ83SaqdhEb62+zU5S0+Ev0DFnC+hgPDNGJTPTQMwnPoJukh5dHqNZcRr/3H+f/0vzD
FwnEAR27uc/wssX+a/TSENSmnuuMAzgfjV2mQjJ6JBrpEetNXg4COnEIUzva6/KJ8T/9lZIPqNUH
k07vPYxSo/wA90f8o8R6MbIN8v96DzvngwXc1fGRhmPMNPC+mwyHnIbkT1ln73+wZDovxcze7Z5L
4vUqvsBtMS/DmZKs0jLA/Kyp/3r38ZK2qlpmv93YadmpSV8s6lawFS05MTjxpHdM8vKHY85Uaxvu
46Em05uF2sQEY/tKrClKWstub/kwtX05CRYYZCT2dSA9XR+Edzu6b51ZoDDjozloS0ZG7BjaFHGa
C7KqwVMOrQzDfYNx3D8YMVJhGAJBEWDVro+8f6QXpD0x6lsa2K57FYwEupcJL+OIuig6ZLHdgYMi
dzZZo2h3jgNAEnux/+Bu95i+7meRy8Gpjc0Ig3oiMijquQ1z8ib0y9kHdLCekiBPyQeP3qBqPFfB
bz4jN3MpiHfvP7Tp/mcNsMj5W9aP1lPRGtp16dit8C2Q3AVz2+SsRvbEpSmwNbTPXFNXcZG9wQb9
/9EiJzKdrzAqS+BNl7SZUz1UmTsSo6Bm127lVgq+RJ0sf8ngoadmFZaWpx6ddX4py2/hD+7aXtgK
C0hJQZEgdS2w78pZ/gSpPiBSJB+6fobFFNegnj2A7zlMciE2V4PInOVOUFo/WqlHoYNbDDFvDAsU
y7QDNvjJrDdNhlUVy7MoQ3FT1U+PFNYWiort+XTa3J7D9+LvcWl9ziJjdYZA6eGzMF5NXQglAEh3
PxgWyxW2ix/tVd+hdH9q7yGQ+0eLcIohsle4IexWnGJnZ/1qcP96wplcvK4EMDcUyDFCiUIdtZAw
TpAuG9Afp0cOU+pRMS7Mr1YRs+cevgc9233N9lBoO6n+wf2PvPofp5GptwWAYeQfjWKo4/nD5qXU
YpNX8wRtoP+czGb/By1gGqjQNmMlYN1j+aM8wjsRjHqcXfWKRsrPajRwCyUHtCpqywNWdmuJmjhH
AGvMKid5MTxaoPyUZP2xsD4XDeViQEP17Y7Yj8bTR+f5lC4ZS4gRvd7k2t0ST4Iv1siE6Q0ygF7d
r+3JMYRPhVYz0e+vo+2JEKRpbkw2AkjvsiAyxrsWnE1klXirff6zhx1Wt99JMocloSTsRRJNgK5g
N/LcPqP97DL1zVvvyFol4PdC0m6k+v1nC8fLzFLywObdNBIsU3dWfCPEiUl2Lkk7X4j9+OyeChlb
61TduHpEkhmnMqlEa57ZAlMEks+YVmjBe/14qJaN8FXK/J7WG9pY0Bn6gz4Fzlo3zvTZZtawO/dP
AUlP4ls0+OzgOKMSNsaeP2YeEFqJlCl43Brh9W5UR0sTV/QooiV+x/N59XhAItyPjZxVs4+JlpsI
dM6Gfxag3Vi1E192kEChp8elCGRNFAhyhZaf5gkWfzjGA/s3g6vHXoi9Kbxi3C2mm5UmSlb+yljh
dRONQDR7UNllLtzHDSfhs2l3VsrgvQ4cwbXpT3pxCZYZt9dgDnnLDZTY4VHezs1i7FT5lIUjtBeE
aKhumxgdBzgivvHpVOIYBSVAtZM3c+LhprjvHa+oD48T2WvfgZqtb9UmDwoByJEW4UM39Z1RnnwK
pXNX9yxa+btbmZ2r0yNoCmp3ZoAdpowbFThbQ0HoYElJtor+pBRw+pld8bcSUfJFe9tW0oGfpe/u
Gy3VTJycNyh2/Au64RhWd/XXYmpl0H6M3JZHdoNAORxJRpijlLSE+OY5uTwxlWt4ePi7am4MLQuo
jWCOltOrfkcmFEzmjUxIfEdqnDXfBLK1JYPB5H/SB5QxvGCFWBDI2zOBzx1RkOm9lhiUUPIbFBcw
3QeIf6LF1D2IxOnqT+u7kAJ1WBlqmc6befadVzuMMoUihmZIalkMzMVYeUILLBWOQMeeqC6RJKDh
0CYp6BCmBVqsalaw4UWS+5xonKkHehlCOKH0EesQc5uL8TXGg5LbHDI2Y6WXmTAx7RDiJhcnTweI
+DV0PmImY2pflc9xoZjuO5QCcUiA/opMBuZdD+QU2Jy5In/DWkkLckAFUraS8Sj5tSdGJO/tls+A
vwOTzjwYwtlS9AxJQgtpXPpAHpjAuOHui5mf6pL/YDU9uFMG9Ugr+EkdFm6xTahXKUDaND3DkZRS
yJzaVCl/cdkxDOQHvupb77zn2BBCxYK0NMFCK/g0sl8DaizOdWSM/Cbjwl0tB9tEzhtvjqM7osD4
Ab61qINzlqyR2zf6MXBXQR0Y9hdZjMr2qXiR5nLqB63jOKTFcbmde2bt3K8uTBbB4e870Q2u5oy+
aX5qMfeG966/DRpI/fGsw0lzODfiyfuIYzo/H5gbt7kFLD/eTrM8wnewoHDmTPzCrTPW8LoKzM18
MWr+u0v5JAxriqhlu3xHlS1+MMctcivO1Mrm2PtdPVEfnKmZ21vwQha4l3SVxLyyCXgMsblAqc2d
5cIsbhUGJ0HHeLoOdIiUNe/joIwX5Vy79xGfX+mEk1LI4FZVGEWZ/aB4fWjDTgxKfx//Ie7CA9FW
zb6IWeO8qfBcEE6H6SdZNugfY2hr4hHazzTI53DU9bb/K4aoxL2Rh6Fn3ACQJS8YMGz7f/so47b9
8Bw9QrmMqM9pqWq195biY2b5737iP9NVYeTpgryk5DeeaQ4GCIPze6R4BEv1NAADMI1Lb0OoXPVU
3Da4kyUN7kq6cHqNd4M3xHCfpucBBiRantrCETFFWNwWM8HYbwEeCtpgRFPmqIuGT5XRV1D3VQ1D
QKzljqqeBh04fuEAbbZH5cWnDQ/bPFDIhJrNo95cuo1lvayoS4btLPV/Oz/yF0a/zYx2dODrPLQJ
rsn9ELVCWHZLSrmoBneYUWtiUJTym0SMUdq6tTGMRmBQVplzh8gmTF6DiiDDu78rDdkFg9kKXTh8
igZMFaNv7hEIhaH29sUj76ZHWigmXYHQm2Y11qgJXTPGBIesWNCpEPwN2azMI2fRVftYr5bOt7x/
QFBb+4y+bQ3MMht/QI/wXylkvlJnEwm3VIoy5GfPgKPdM4SEie54D3vERqCn1xfCwaCgBOk2lnKz
Z1MjEycFkQupPGpbOSPJFk9c4DTGxW/KS3J6rX9R2FFZYI2SMmYK8If9gZDszsPAfjsOkwYdflAT
wQATdPwqeMYnjRsjc5xuCIzFJ+/kOphL73dtd1wEccpoDwiekHknbiG/XLIZHCTyr3dRkhQa4fJz
dpdEkjxZPiuq5dtS2hebg7UZcm4xDMO1yDKcjwnOQ89zEhVvTWlb/FPHvVXAorTjVVHJyXbHyWFx
t5YmBopAq4DFD+UX3yVLkpju6wHBxr4mnI7NpNhkDPjdH0G5z5aonpAFGANPNpcvufWF/EH4Ivtq
axezqa8P5abddCcpb2MYHINQXUqPzYGrzBsNppg6UZS0MYDMs5vqkx7sr+x4Dt0NS8Yhuo3Fy8vn
w/Pgwv/lvSNqLdZI9+u8mEFeSva9gD0BuB2zDpYdrKnl1GoeqgYfP4lLKJXAlfJgPEGjH6ofXdZP
zfQEyLGEnxc0x4uLXfcS2VNEV6m9uszpcFQaYgaDzvBfN8jNYhVOVrDctFT9SPPyfzGxZuyWm+0/
pt0hfQ3kJ5Erm57RwnUNtRUnxZ1xo+QcArE2sF1sSZ2yQSheogzAb2lxOvDqocDYJBKNVuEwiiLl
as3LglKirDV2KOu23koszpFwVv2KiGMc+fJdceO4Wa+ryuorDYvAxBiqt4zF0wp8/Ajn5BZ9YVHn
ROKtI/NObjmCBlpgQ5hCYWu+r3gfQx5VWaINs6Z2tD9r8czc2CPh9EktqjWE0fJMue3byXyEhbVK
FEQuHnZ/1JU6P1YvTql1YHMuWoWWyL8J1MGLAWLajDiBD/9b51IEV6/KzpVpj9zH12x7zzuXkI7+
s2oW8N5ICKOl8Pcs6y+kOOOlGtKiAkpJ6JktiPJMFEfRv5LWW58blROm705BjGrbWA47fkcC9meF
00X9v/9rUXChxkTjy8sYJpAsI9WMQ5HZtKI5+56XQ4nmbm/srNtEUnwJziIjEo7D+zBIkmEZRGNg
jKFH9hfjD3YOeMYgOMF1RDbguLs+J4/Z6peDRgw0drLxpsv3cqBwieetCJsn5r0qqUwWHvgZoqIT
PR0/YlUGiOE2293v2Yt33t3z9lNadaZHUQks82BSj970mG7nHcTd9iqetXSC2I9JAAVVFhTFAWkT
4O3Se9KwuSGLRTMD1e0d4s6sQHUDl88TkEf5SWYrJcdKpZ6QCiIxH0xJ6kwwv5mepNXAKTYsEE+r
0wbijlBoFDOElOA/KVHIdDwjm+XbkFdO1SNZa0AYyoGZ991d5lkA43oVRf17q2tERLHK7bQ7aDIl
pDw98NNMimcFqfW+vGvNtPqqm7cI0L/FZVxXOg3mcvDCfxU1R/OcD8vDRTWTBS9W/BH9aU+L0Psd
dwNk5OHLwgOxsQyLJB/DPqmNuGt2m2L0zVnSz5cn0w5jsRtA1sJcWmx7vHZC3E2aJ20DfiC4GKJD
WG01ZaXNIPjUC0Q5lkM2p+m5EfDNosTqgBr6ESGkpON2bLSfRmDtPowNaReP4ViOg6jgdXkMF54/
ZkPda5GRTt6ZQf0yTBKPfEmbA/bD2p13Yo0nIOD6UU8LW/uUEMxmezQ+X+HlUxrPu2aGJc7DfZkM
eQJAXmPga4fK46UPjrlNAiVCcEOj3UmaWww2uaK4fHTA++o/s9TqGTvwRMSj9elpPhQ5O/Jqh2Jg
Ssgp8W9dSvbxtZMBRD64wPuQoIJ55pjj5wUfiThHOauPe4oeFYEyxMxg95NOYC2KFxJo8KX2v4TA
hh9GjBfY7TF8ReA6wtUEuWVmYXJVW0Z+yhRiCpOvNiCbtTGEPfSLUJXQp499B+GGMpGehJDsQOOR
0NDrwuMmLzmZOihQvIUdFon+DTd7EnDEGRZy4K6iHhNLmrTKwN2WXImuL/e3Dy2S4s0DWM8+T39+
YOriv3GrC87k4F8sDVbPygbCUs1FQFpifRQYozvm0P+cwt9n9IkkrHwlxP6RpOrcE66kHtLQi4S7
xaAvFC/PIglHKVYFLojcUmnmb1oiszGAJm5SaGOPWC4/9JMVJl1PjRPwqssLBKCMZ8mGizdSu8/a
8VlV30ABhrz0HigkFI+ByBBDMWhUl1KCTp/50Bk+DJQ/1P+B8ah26x2XopFtf7iSYONCUA4Jifqq
+1pALY1lYTQlhRQl41xpl45IrjvduR6fR5L35Z9sxCEBuhIVO4FcQhfjTJmXYPzsKlF2hmTPAHR3
6DP2XShgPN73Xtp9NjKrxe22jLzTEjWl0znbhxHB94NsyJLDM01WLBlyO2djMBAQvo9n9eQRaIHM
NugpSJgNIj+5VDBvw1TYylAwrtb0iBJ89sEXmoyQQ/NdfQ3SY09MSX6a8pXtLoMvqN6zVFXnMeyx
Qehpz7ARhJF4gYdBnuUHEaK3S6qDbueVt0NOJZfV7BIz+rTXOJvU4Qi2NSRmSAuoDB1lUZfAvID+
1i5MSRJwZI0Tx0WaTPz1pIThgAGCID6ni8WlnJSjSgKeR0HKmcZYMndbMPRsW4+FUa8929v9/4T0
ZLB8NMUO1fse5GPfPYtOjDtFYTE0weKslsVVE00sg0T5qCou/wJx32DN6GwLGkZn/OeCqoV8UK77
Rfbq8wASX9oX2UK2yW5wHSt9HnNkgIQhwYPpYcuxgtfIrtm/5/xGLItxcfLBVKtdGAv7vB/HhJhX
62Sj87UjCLdkfwpL4LbG8IIdcYqKTyOEZNduJVh5g3RpHKyMuE6JzFg5FKS4aTWzdvyAfShBDzyk
zGnAA2p2pCItETmCgNtTk1CCkAz+gXf/SZe+6HIGLmbFM6wuzO3WqD0Vnom7oIaznzXQ0ihFNvFQ
WILPlRqnXOgNKVU0bLq15X4GYeKLg7Nszx8JhCCtOZ5KgigC9vehjjVSOqAMF3zV3aARhD4SlkjJ
YJvgk5enL9o0C1+MkcmAzmxRuQU9kKJuuWRE+38dmo2UHhAKv9gdn1wF4ybffEnC/iiEH5ogNMqR
5NBb1dllJVotj+XGl30tx7+U6MyavKXS7IIDkM3pDq0rRbjWPY2OyFWe0HDImk0MAoXc4bVG/ld5
QDPVhSCxkBJ/Z/xyvwXhxvKoQqo/y6MfVPrm3vcAXZ2nWfGIhqNaFWhZx7V/8VgjedTnJjYyZAkB
RVfvjg9SaSl3rrugMuFxAJV045YUBwxW+uet8HP3MD7jDeNFeI27Nl+9WBWUF/06ZIraSyl/kuOM
sMAkCu1oeX/+vPxG7WRfV6S8HrPkvJyanMHQ4nkRego25fpcUlx3VLTq00zoUGPeFSNXQ7esBl/W
4PrWMGsHPdA/H8GeduytX7x8tBrGgkNgGw3dffxJWLTbZedD8GlE/KS8EoN8AaOQ8gVV0OSbfbFD
8QGXagI3q3mj7CTegQx25bTsDQ+/iZI5MORAcoUcwi2noceZGeQcPhGJ+/0PyW3WVpUBAKMSK0lj
TVZTjU2q5PNSblj/KOct7TKrUhuk4bHs9QZtgdlMlsbpwOD1wPhe8XLPMu1xW7viYx3KLJvSmjQI
oGyKJk6Zq6Gk5Rybimg2G7TVBeBDnvvbZQUebwXqDjNOp6k3O+0fHdbjVWvfl8QAtO+/CBPFr6wq
1V5MspvDxPF5+wQy4L6z5EFK1SMwczUVveV+4ZSFcpNrOPfp+v66ZgDge8FjRmHYIsZCuHYCd7Cc
TuVHt6Voaq7q21Ty8oZ8Gt9yvl+D2cgRaSoyq2II9f1ma/Rilu8DbTPWCZbOgzXU48YB2mp0LGP+
XlliDfapAfrW2a7qgAVL3sIae6NWPaDKImZh3p1yJO3Euva5krB8mduWku6vyPXbHPWlcYFY/J0Y
gLRv9jaKoX1jdhzNQNOaKuIzLV+mDBRrKM/9CIcRWZwcI/pXN4q974d/AfmwQG2jIGJP3fqvSg+Z
bVSBIexcRqicx/AEU+IrnIPLVduO18l4kYfwve4ouAu7pd5ZFrx27rrqaBUcU2kMoN2ZEjq7dGr+
5WDw+9y5F33fVIuK24aCYIhQvq5nbm7iKJ4X8nsagG/rNsBzFcw5cQQKsQ32AIdsfbsbjVYbmBAE
bfnJWXIMaudiFvruCyo7Mf5XFXvLMui0+RCc7eWhwhNqSYusTefQuICXZmcf7zUcwQnh/+/E8CXb
ETI/DaGcqbwhQei0To9M+3ooVaf6V8ImxcEqW8ainx/yCWWd76ckRWewBcJQSh9kwuVz6eZt7dWg
8IW69jFSydQxO/LiQE8g7jU1c6PD8A1wRRl/WU1mqhAcTz/TkbUJkPpJiszOnUIlBmPljtsTHZr4
xQslDvGnizoWs160qFmGXt6/h54/GHSn2XaL30CR+UvRfrvawm6MPb4X17b5Stgw9y9QUlqm0PEO
owEDSbXWRYNdhWgnpoPUw+W2C2F8jyl/9wNxugtXgJ3JyODsYfOCY5llMq/JwDUMzrrN8t8z69wQ
heFeJLCSeADiTP5t1PKtMA6gs3YDZr1i9WKPxdwwlky6TlaCWmEbuVe3JKUb7AgS+BT2gyX/LgEM
ekMky1ql+H/U1nuBi7Gp0wZsy4pOTZ7aCUsb8g7hQSYJW/Sh0Tt1PvYa9UlIr/lS7CWhzp7TWpRN
yEQEAWgZV4QxgwrL7Qar6Y24XsEQDdnofNZ2gjWgAP69VDPFzDv1Mm+uMvHP13XNNNbVFNhF831w
d4T4PI9uIYhRAkKAocHP72yRt6krf4vgfLWWJM1rUQ6tJVlzGXSu5nlf21tQw+fqqtyFLqJRxcCA
8ClMX29yHj7isBv4J0HqzRXwwAXLuHIo1PxbN6KGVfxeltqSQHEPWgPef5hreW1mYf6vsTerIdOu
A68Rrk1hyG5IYKVgcIKwHTiW/sYjsvjY2xNyK8exXS9fRVZCYWVPfLiah2TisOQV6Jl9m7KXA4NZ
0g1Z2OH8Y0H+1QpqrM6cEb6FT2mf4pJIwXpk2u2tFYrvivioeRmszqnrW5apKOqRveYYU7dLt/31
fnOF4660i9ZoDTr8z3ThOBEehphcIcd35fpi+E5Kmo3DAaed5yJvn4HdkW1PQUZjfrUdT+zhxqy4
kQpgMVFl8z+r5ox62k5eI+mqX4GmgdubesIcHFfkwB1HnWU2V5UTDQYk96Xc3NCuvFym2rRCeeGU
WTYy1XV0ga5kMk/vG6oMYFgOLtKa4pMDNzf3sSnsU/1ZOp59MjZe5lwp9GwoXek98CqWM0rzuSJL
stcQVxg/gY7P6jZIMid5RXz5/If7MQ2mhaMP8T5G/ZlhLvFOrZD61geOz6h+qrhFnXJaRvQs6CHD
GnxNu5EF1xD7k3JDQ6J8i1z8PEWI6zs2CVRNAWfw7akjh3oiFqNPg0JIKGNkHU4HPS8ls1DxkEgR
Bimur+nYwjEvp6lykQQzykt6ugi0eJEBM9hL72GIXj3h1nf5DdtjYlPJ25/MNQGQz7wkC/9Y5ws3
Q6cAxLnpsHC7nq929/mbxOZnwdwVT8xdDeI+LljYZ+9rqJL0U8cpm6k9E7BGsRrxAj98TtuIIjW5
kXZI4i5y5E3XaIg6wJ2dIhXN+3noc/iVbsyXTVkz9x3msuE7jmm0efLNUaDyFTf0Cf2BM+Lux3+m
YpVwqWT21bOp5YnTF8OYRMGe/209+SLVDrDABBCP52JLPTh5Zqt01m9zE39F3vxv1dC77DEdyRAb
VXoPUuxw2w4CU/wnTAkC/Oa0xYmVHdn/w6VE/VTu8ZsVM66avumFMJ1MAJI+CJmRPxGiCxz7SJ8J
Y8uh1EZbA0fWdMe3GEsUea2FsA2V4mPzOj0meQSyZE8kqi6Nbq7gWyh0vB3Kn3SMYEV0eH3Z8FBz
Srhi+OEncIrwaXQlDyebpGefw1zgohsSeql+VqKFeHaOw4kaMT+z4NN2XStMtGTgsjnGozmRFhbI
YQYXpePUu9R5ZoQZnZ0MNq2M+jEsrUgm+PJjL66Wz+gMIL7faXRX5/hMOmoSmlJCVUaiHord5QRC
3v9B+c1LZKTOoBbS7gJ42hqc8+sFHxCBopAwRxDaMHtzeEHBaC4OwGQ5RmqnlDa9nDBeKUWsFrgr
r68pjAtAKBxf1I9y88XJPYWGDLhwwb5gFyB30qmtU/LPGl98F+19q/WC20BKAju9hC8vGiZd5lnw
cwY1lG7noFv1B5gFUEn1ofT/phODrZJWuFCN7qnnnrBb6CuKGANRb6maVoDpb0iWzKUvqC7GTaBW
1XR8ZA/WHFc5RJTLq+6zGllhhjwgj+84brdH6PugqigA3/hbZA9WnUxuEGGyLkOjEIY0AOBXR6Wl
gwKxE9vvQ7ZY+tPiV6KL2Ft+CTXNjTgy0h9G14xrc1PVqqGq+notjOfIpYPNBRDhNFEjhu5e+CBV
Hw/clFujco4uKidJIoSXTwrZ5u2P+S16aEcrs6tolt2F/15qPd4X69Pfj1kwbdWMAoKZxVUsnt2F
ON9PP3jb2bfwxEmyYXHNonv7JEVC25svYOUSJ49kZjILIshs4Um+Ditno47dzUA1bxolCC7ZGGJN
+80BJR4unxjt//LZoG6Sw52y/cgBJ1Mo5Pb76vn9A43XBTjwINUS1LpKMMNFSYlgH50Gp8ZHjBAq
U4mZqBR08DZ8tp5PCycz7CI6CqCm7Om8lC2lfvPdyVnsdcycj+TwWdq+2WENZafLAE2eKnVJKGt8
WpurcGF9OdlkZpTWexoD6yzWrCDifLbtGEOLD1blkEcy7uNC2mcirAqoD/TjXpl9Au46P9VwWO4T
AoqHLbjHNPh5exEOTrNeOw5mSE4L8DbhNh3udFLZjPSUKM6pj4rG+UoItezv1VVddIt0j0gcOoAc
5XfIYwzKMZwa1Eqr+U+cfpa+ldx1+x89bhqDX5m9ye0eHDb97AmcfrzAWq4tFdg5V1KVy3y9X27N
ond6qpPA1nDQTzN1rGG+6H1mLx64aobFIlz1KVpTE8jxOkbmJD2MVvCsW8rwU1oCd2fNALxVDxt+
MSQDG+qHeY9dJqHEQi6jJyeBhws9GPTrEiBDuvCXVei83fb0WTyilQ1Sb7ADMuiBNYPyR6pCZprA
CH/hj4dca5JvIEbXQ25xE5x1odHIyFldLStnqXALbOXI53Wolj5ZNfuCxca29i6GiETB/XP7LTU5
u3nwtsl8CKZKmxH6RLMU/Uqem6yC24cj61XhbVmMFsP0Miyi+RNkQeZq/OibIJqEqGg7MmMVGm/c
7Sxq2kKLxuj2O9MB6FSE5ogqMqsPXVo7yk30kpnYorUfMLeL9eMCVMnuA5DytuW9ysbTOmmei9od
QhwIzl1dD8AUIODvKRGSTP6x+cAJQn1AfyqHcITwpHdaJTrrCNrgOp1l7GfPed5H81xsWfFR31+0
Qs2oW86xR4E11j5gN9x/q+oLjUZJHFzFTvLMolAj+g/2lxARCPFUgZjHtD7FTNfdcrxJUyVcFeAP
deCGb2+sASVBipKjf/obmn7Rkz1SsPoOeeONCZuqgTs+jXvGTOFn5CLu3S6awhypefc8oG3W/Sh2
xkl2iUIYVKHHxuQAl2G+9wO8Sk5xScWXWhHANVVb8JFIhKAlCqAhwMNqPN3fqCM+MD9eGxop5Yht
ezFVlU8wZfMFV8ulwHoJ/YIHsxtXPJOO01kF/Z1JTxsNdTxer3sLbsr1U3LV5USUFJm/iHgdpG48
6JeDiy67gSkiWBvdi5aSuaSlAECj2Oey7KPhOf5+485533v0wBh8I9XnbzIylXWyyjZCLsON1r2m
Iydl16+0VfjVqUxdNzP4jVhOqe014cj38E3fmhPdLTGSeNbFOJmwvnf6JYEmOqiOwiKt/cWXJBEG
lLfTrEEsOXmGOvV3PWu6hUcPX+mn35C1AH8cjU0xCk1xcad80sYyJEjSDLvVPvG+yewi1nJWZ7NR
0TiVP5NqhOl7WHVtytb6gDrDqRdQFISd4LGIiu+7JXeTtw5E9K2VTeCw8SKdm6Z2atEcOzNsbHdK
quKLDHhutOCFDRKxIaDSUx0Fc+DgDWbupyGTtZLAVcODbOfvtMCww9EqyqErVp7oVqQwPvR/4Jzu
gNBXpmPFMh3k4EChRk7gmNdPM1F0x1qBx1OV2ceTWfA1s0VhTusbYI4dEP9YDV6hsPKvXt4MoObq
GR6/TfAC3tM99rNu06ZhRTg3aLh+bJ7O7itcyaLxJ125ef8K9bjEtMQZWc4oxlm7iBx93qHjQP5j
e6eoIcUu8M2lKrG5R1yK+yTB1+c1eHXzLDKM8vwCedS5Wn0gmtr4NR0PayeT/7fNJ4jeEtXHDS8j
FM4aaEUyx260sO16/dsiFYXqLsQnK5Ffy0b8OxDLwS1r+GBNTOFyIS8eVN0L+Ao/qaVWg5EmgsWz
EdiylxW4AT5ACqWaRBCaquZy6s5yOUcwA4Mb7UzIRO+xlJU7FWU/lSzeOLtySHrKfPVJf4R+Kcjl
z4AbpMsF0Tc1zoEcGTJ0uCbFzgKUxrC1uEf9dSsrbTRurI4TSpSuuJH/l8U8alB/G1AKZfLJOYF8
/rWUELmAP7yVPH2ZsGR2INsfjwwVtyZ3Vt7sMPvFN2WVMmSmhyBw2eRdEKwerfuNuzDTNW+B7w0C
xek74o+XqXiDWhZ+7ZSQKC5W3cH5U3pwc9jCDrOkjg7nlaR7sw2iBexmnBDcg0yNM+wYQuFFTZbt
ciBULU4M6PcYj1WqanBkhA3Qx3EgsV17t1cTwhActZz9FfVPRe02M1ZDYmkiYpp1J1lH9TKE7wqg
NJM2IU0lLZ5BvAJQJI9C//rfOqceryK+DapJZ5MOwcEj8HIYq7rWFTzWS3aMAmVmhyw22vWvGrkf
FrywRbngQ8eBDPUU3eEgzuyPtD43putMwqCkOf8zhKf75HVTLw/gIup6sOURGP30y4vVIeqKMJce
kXvsI8mWHiYzAFqO9qF9I5RBCv6aRWemVUpe9h399gMca8pjhudItkR/Zhwg9odfSka2CEWhr0as
eWWc2uCAI99iDxQAmAxJy87ImH7kbnKmm7BjoGGhbulf14LC7xCfgsDEqE1bQo9BkFZXC5UfRi5I
LdbRtCKyFvrWSZVm9nxgmpAu8Ek+MiORgAU+nuKyvSeGITcEa3679k8tSJU02FtxHAxt3ClbO7t/
cODCn7ScS6oEC1AqGTEd8d15sYYzASQO2Kmv/I3Sobzg7ke6Y7htImDJYUuXDT+8Q9inVb54wUL7
s6ISrcRHaTOVoYwtu1mB+yAYs9watuz5mHWqRqdAAl7r2f+rkbXnKAiLYTDw6j1EpfyxgfuoqrPm
JPBoXpOfisicMQU/LXkmTPJJTIGQvfbdh2qcW2rvjE2p4Ew5OL1o/6HcgMDA7rEyp8K22f/obmOU
eJYeLx16cddZ585jkarH3nxvw2jgHuv80ixaZXeE1mD31dJyZqfx+gyDOjQ8LFdFj6rY0lEfAY9J
BmMDEuFtHY1hO3UBZPgmaMTHOkJOgASqdDDvKt8cjoTZCm47s5VW42R1Jr334mUKqnxGIvbRWeiL
Sm9n14cKU948JqnqzMiMBJ1MyppeqIerHUWoYoB0l4qbmDVmAxPbXlKu/4omjTpetJNdc1nyJU5C
19T88Ag/Hi+J42qTOjG8Gwa9A49yXdE0phXmu0sBtgvtGPuBLXoa3gF1TDnRPBoMoo4+ZdWCpEvY
uo9HD0/0YQL8RZVZF0h/nXQhu2vBPgawtAu3h4OYiIAB74pY0chePC2Wn13DT5JzEJe6+FcG06gd
3HrcXQ0UUEJ5i7hMV35Xc6q1Xz/pnnvbRmQTcqeZ4cOu8utQJtkjdthSB260QkuJwt/OtGMDtjan
VB6F2umOVx7rx7lX9f5KJdY/cKRWoRrYQ5VCf+l3rc4GPhMfy6MNefTkPEsdgFFOxQzreXX6H0nN
TJ38xPuND8mE+JTS1H4aK2eY31C6S+mNUzwrqUvQM4r5FezvLKZyAJmdKejUFbEzAJOUYNen/9Lc
O1p5X4CMi5oFNYB0uwv+pP8sDm7GtAKw9AYrEWDyEpojB8TxGv+E+8rZNaFpsmhON2LsQr+4IiF0
e1sswVUWFVLCbQxqmLIK3Wy04XbIGXhg57ZeD+pN40EcZsP1H2jLi+iqcb/bo2MXFR0jJRUe8yJ6
MkVVYO7vPzhgEcVCrHr0r9He1v0icsGo2DEWq0P5prccvxRC4Tnb+N1FI2kjMsuJGM+cvswwCSvj
U8vAAbeSwTEw6v8OjFEjXh35CLKvhsiZHu9HsLe4DSR6LHvmFEcNQi4F1z9KZQKngJ9xAtKLmWnx
X8OUI0StePTeGOYP/qkkb2jOrCD7Ng7LsF8ASKSNKCz4uo8ZI0bs+i8yMCM03eb37MioCNdjyZ+v
WZmdFuZUaE1lRseEQpYKVaZ/XnibXxWnr/5AoeQmMMym42qEboXRGSBIECr9/1vQT5E7SgRqao89
KXwgkPq1UKB7D1TAtZH23UYgrEB0OlqHHk0p6HCQb9YoRc+/0LFSjSAbTArQ07xpb9I4BxFwsqHl
MFKUkYQQ2jGODPRmupeSlruOUS006/2ryawfHyAga2l3tntvKVV9WoW6YciIZyquUpjFRpjuzzow
+wVaeax+3Cfxskwj2R91gk84cyPAnXzyjdsMXoyLHLwMpaqMzXqkrUZkRCJz66g5D7+uh6qOGoov
fWghVDZpSZCIB5pB75RI/NaQgv/gXnzWKap3KQ42taBIYzkA3X1uRM+yr7lUsdlYvZOQl6GyelWd
qf2BdCfNOos+MwBugEflEHSn1cmvu+FmadVzIDLTgecSPRtLjek40WUlmxI2FB3C6NjyBDGsILZY
ZErY6CGRIDTMNyIh7RAqsLO2NI3eYXcaCrIf0ePSxcxlQUl0IgSrlTBLUDN0360EA1cjKhq6Rvzr
q0kW9NUNbo7vSF9StJH2OxxwNDdt40eGhCz5VdWrAc5TBVOL/bF5ZybxGIcRW3DHnCMpjLI/ebgp
x6wB7p3qzL5vBcS9WFVdYlyC4R1sJU1aw/4T3JrRXGDjPe/0MmebnbSKsnCubIGtVUo8/nPcbq6Z
MXf1z+MESs65zMoxdtJAXM4JzQ8XDPAm8MT5NjAZMPaFVXAgnZn5ivL+KSRepwLJJFIZjEP+oxRs
NJcq+e3Ps7xqen1kdfNmk0kPJ8oKP830+trKVa+J3yQMrri6PV3Me9uAPQsc6aFpMMVG/Ft4eH8i
kaGmqgTxgl+tfJcbzYnsRvp3KZ+XJ394n0OBh0dpYhdLE18upPkZ8f7grffyIoYdDBG9bXgzqhRX
FexHrziKVJAr2nTHxhxZtbyu2LPDHZnjKj8o68Sfppx+ZYdS8Er5iI4s/Tz4FhqiinOS+eB1W+tT
3maV2PIOKUXR3g4TKnNXne6dNgpKCgR68eyJc93nkFGwJgOfBWJhNT6WxI4kt9oYuEhb8zxLWcmz
0LqPohe7IOc24ZoyedG6zr81QyrZ9C/2u0QwwK0tDPFC1RFC+PWvtUqoSXodrR6E2VELvHl6oX+8
yJ2CtdhD3LdvXCeMNjSV6P9V8h65Nz+BnpY0NOIhcZZWGSRHdDd/aFIVPfLXjgs+0DnUUcrr/lmk
RHB6xdJo7pXG7Q7muWhwFqDD7UzvqwVrOwYjfbjVlrtaDNhjiQTUGkPY1j8YnOGtxGq3cxEPnMdK
QOTo/7ccOiMBPiXQY2KSZ3Kv9eBDHdo7kY+Ya/u847ta6e/r7ltPrNyOQFjkr9SN2r1oCuioRPl1
XDZhCjHAu3XCzfhokIVPQSc+OQwsCHat7/MgM9ZdQTNQGWO/FtzO5NkDdcuPUoMrhG16Qj/2Nris
Hfc9Yfov4XkxGwvE0pNrODddAxtCU+UvsjutY3nt6fLnveDd5zfpSEVe3rGUZvqCygAENDurRcSU
deQfv5SI++HZnABsY5EPglKoP2efaqNVaHDBGq/IXWnsvSatUEv+j2E6jOKx2471epqGagIgLmLb
cUBPHZwAKxN9FDeIm77m7nZQVpWUt27+bfLCFXaj3aAQFBKlJXUaRcrjX8VvdJ1blU2Ng7nyVB73
2Vg+ms1DrgQzOiuFHDL7aIa4WgBdIgf4c4Fa3aamegaI5kTpkQCkuT4gOZkRdBr2rYMvymUV3BxA
vXSHYNnJQVbk4CplivEp2vdrP79TAXCeW0i+WPIxEaNd2hWGpP79sohOlxJ8JuoQvurmp/UWYafz
0op7+GvnESoHzdSL19sGHJbdwq7tNC2lv3XQDyVO5Y/dgpi9DhBG1ETz970CLeGWYCQi8HoqCO5H
6vHE1c8n+sOWTGegpvHdiHkxe1SLUyyMwSDKe/jPD5Nw073dWlog7u8FBEXIrxvfRxjGTijtbPC1
hPyofHt1q7Pr7nFPnDxRmxT8lhPPLmncWsoTC+wMFYPjVuC+TRstVnEZ/YXSxzwDWV/iCT3NNGen
MU/FV5TfaH3FXsUtiuXrDAqWLJhiePLIVNYTS4dvCEubjKq1pR3X7BIBicvSJZCXNDnJEVEm+r81
tqJ705OkOQNUyo5mLczySne7xkn4oIFnHfAkLoW/YdYTIKzR1hUM8k+ZwIf/fEOHY1LJoxUqUtfw
mo2dJgAdGAB1DXh41GrxWUK9OIbpAimP+YKL+CLoRVCrZR+Nz2iQSXDXJw12GFTdl3wQ+EjKrIsb
W856tVUbghEo3c6kxD57FRu0xnTitXs/YEj3kQigmelizGpQzHp2im7sqGko1Bondp9kWnS0PEYC
gIjufydnbB56evAaIVIFvEnJ+zEfn1A3HyaSba6ixxLUrljb1PtCw/infQo9ZvZhNcTq0/hFdUCL
YGEPJJl5Woq/8ludctcMWT5wsWsw9flcIcGkmenkn1rd6x1EpuuGLYvN4EvblXrTmfJ0J1Vn97Sa
7aUagyM8a9h20p59Z0yzxQ7JKR1db80qgCltDboBzOPrfrwvyzWeZ8SGipRxgZFFZRZRipQNxILy
/5IMwGFHWdv8ZW0IyvFQUcavHMZ+QRqwNj3+ncEtuA92O2MTHPvjr3qC8YBLh2G5Sb1NXW2MsC8Z
6wk9FWP6mbess5oF9NcYONkm9ZGU1S4DKv8hlkGqD9kkhyifC64ZpafJ9fzeDI2YO/5xmvPiupXb
Y9WbWnESgvz+htFflCOKTBZAW5EiUyzuErbk75pCdAvIiDXdCNSDmM/tWuNqhUjodqSjHIku1K5M
Ir/iOfS79sdApojM66uXZ5XY/pvTOVRlKbrl/iMJgUxW/WUA9/eicsyZ0v2M0NR7YLLLby9PDSqb
owwUhhyZKm67Y5ksBzRcVdhhD79k4jyIAEQLdJHK1vRxAO2/zJwoPj1f3w0BWFr9Y3TstfjbpGD3
XtcXhx/qMAeuTszJXwmGJxh9rzEW5LiYZHKg09Viuaqa9qNMyotR6dv2i5v7Mb2xLAkKSHz8vVwp
Fzob6dGmILQKmBC88o/4DiXJQp8amFvBqqWjq71DQHXe3S6usXGQvLRIXzvheIOTLhYwQvPKqzaJ
B7hR1Zq3mzuT+45lH1aHnj9+FuClA5inu5stzth8TFXAgLLq65XP3bn+pj7hPa1ShHZiuoP/2NKD
YM+fIt60owVZQ6AVOLBD1j0RdL8vcknPVXnLvevC2OG1eA7wvyzVdzGhxL8uav+/TiGiQhSzOqan
qj3CzZ8W2AJJMsmOS3sop7v7hF/HYg0Gw6OwjjpRK1rFktpPC3ixpZ/xXsVaQSf91P23GztzprZ8
hl1MQwAsO+qbE4yS4vxTRDOe9nj0W7gOfuEbsAZ7tZPmx0K7kv3tOW4OEX1x/pTGH095VyDzlEvx
Sn+L+gr8kYv0rDcbZnzhj8IysvPrvi2l2Lf3t4PDaRCHL+lhNhg07egllgUVJcsRz96hukhB3+3N
Tj+BnpinE7D+E8nNldF4liBp5tzjckB+dl/v70U+fWFgAzyzFet67SQSQDHVPR5KRlc6dtViEU28
zdaJWCK2Ovyci+Gd4jK9O7bsQEW9/qBuoF1xZFnkaqS6gLU1m4+UuOMI/MtpvN6r87CRpHcuR62c
4SevaCx9pQez++mTasMia2G/2zbuzyPsMTHUwYF4py49lcySNWBKIKvdnLRY5MfGVSyAZQrotZDv
QwYe2wmHjFwVanc6nlMdMcjYmCOhD8C8dXDat9C3IaSg0R61/jwPugsrFPNMlOBgfqliTi2/vSdz
FCLuEaPCgmA5sCS0OwF9J9GyapxYbrqUT715uGNQT42k844s2DR2BEZ/G/livv+xFlbrERS1cYH7
Cc7g+Z3mLhhzdZb9WBIgBlcgr0S8XChBie/GQ2ck5RmzNZdvQSlkg4zbDLPL9llu7i6lQTMUh+Qn
MHW+PVqDv/lILnxFN0b7wpGYwI31QwZFMU5DG9+7NFRBerlGSclnNEtXVtRcaMWCo/I28E5vt6yp
PjRpt2IgJ8z4dEfGhLyfF7b4yUdXZnQPRUrYRDL6lDwOO3+EiNrxrwwj4wJUACi19rbcGstc4/PX
opfdekM8LlUCgvvxwp/+baYL744QKXYGMWJt6Rt5OvF9XVUbsoBxOpA01qSOJ/V3Bo7+TmTAfR82
XGSmZp8hYw5HUk3X8ggtiomOMcPLvNzxwtp52FHBrJZDu07RPQ0cToUyCW3GgJY4bdbuWSTgZb/M
fSTyu0WZMc9idinJjI/kEpo7lt0plS/9EIBDr1YovVOCAokVtZmkocQzuco2utpvYShkc8PMCU8c
aq7z6ir4kHF/aa8k4pfb/tvDrfreBUNQQkuHLhK7TbF+7+aJbbR5uLPC4WdUwC24tUk7pf6J1h0P
3BtIoXaJi22vZ0QJd/gzsxkUlx2kFVBrEZ2j8cMzTWLL90zvAaHXCCdCD01STP0VoBZ633XK9MQT
UtsB0KfZp2rZBq3YAZYsFSYhHQtK7JOAbyB91qa+h8+z0khY8w+R9M9KmVwelz5ECsCoPvQzsp6D
iNJp8Bt6+EuO08K6NWtGr70i0oMPE6HZJxx2R+rPRSSTT7fHRlVeAMQyz6HJgtgdLQijzOLNcvVh
QGEy+aJqgFYpWJD9raZG7ib3EINZF5sxzcjEKZtYy1Wi6L7alwzgyY3VKZXn6kE7B5Z88BpU0Yyy
J1VOoMkrWJ4h8pVp/ij26cT1I2XPMGRPqEYjp294HLjVgcKd5kLM+OT/IN0J8ZTiXqRabP45KtJj
06Mp2m374dDOSgwK8ajFOLGYXl94gkRRWuQ/s0vMnSTaddQd9f9o7sXEDjsI4WGfsavszW1vbqLD
QBJTreJxMW1Fpl3v4+TBFCxPDzD4M5jg2vZPJRX/0Ql1ThPs9NvLE9KCrG+N3wjoRTyTyTNkZ2ov
fyIyoW84SZNCwhnwLBMqNqZ9pmDtArOc3r+dZdHb84b0b/L366UPAiH2T8sqjKdN7dBL5aS2idkY
+iYFaFpfJGii03d7a5NcHu39dBjBJJLWAo3t3WWL9Ylvgfxqd2da82/U3HLgXTReKh1+ewC8aF7W
0ThkjvCaYo+Y+mIHTu7OsYNTSpnGUOFFyUJ2HRG/a/BwAGhTi6uFPIHh509CppnqiGDxn4TCgG/g
5ChYCWVIVXkkIpKEBWpkgXD33CLTcfAH/Sn0b/wzpRAwGxxhHIsQ7waiNX7fjshf3oA3EdnsIMMA
7a7zwj2Nr+zd3FMPyKVq/y0TYxtWRK23P8UpHnb9H6oOgeajobwZSYxmkXYUhztNpkYtKdxngO3W
7oWMYfa5HVr0LDUnl3hqqhWcmg4K3gmOT309EGnYSOUuHxDVTg1GpWFvXtGzBN53DOVhJTfxIqlz
TFQJuDdLcpZkSC8i+n94j5gCNGygePf8J6DvdxwhQPhaT+Ne6KGYkaIX/A73lvEC2SfeRWW8vkw+
sBCi/ohPzDavT4SqUt/IbUV3OTYvOQfUtLQ4FNfyH+F92OJvzmBL9cK4v7zH8mLvW/c14D9JGS/l
xyt2bG6Fh4cUQXFb2Yda/2KeeqH8YGmHQh6p14i4XnfxKps1NNTsJLityPPBsnzqf8qgZ8AVi0n3
t3fI3WwR0Srxjg1YjqmBmRIdp8Q5so/d3igxYpsecawnrWiqeP4EYsRSRTJKzR1GM8BxpFYWccc0
2O+CdQ1QtfWIAQZ0NKAj2r/YcTy0RL2TUZXPWDKJM3bE+T3ti9sGah9+/ruGtnKiI0e52CuAawcE
H8M/0VDo2S4xzfc5517LmU57NI6etN+U35xPliVosM6unZ1D0RkOpnyJXTJkmwJtz/5/8sYz3XEI
R2Zd0BW5RhFANGqjWyQPWLJCWqte36af87ZYwfs3E4Na0HREkeBdojmdUHTh9DMoORdOc4lTDxQi
cPKDN9BGwCIrGxXLEfk7fpa6Gy0V3ZWQWQGoTIFJpaXKvkUndKCe1Jx+sJmx8vqFTJb1G6y5800g
VYGznCYnFqQMxh0xKuZEvYMVoa4lcWnkUJJd/KzC+Uq3rZ8UiGnO30QoIPMsZfzuSX1pR2uVuYgI
6/XZfX1DgFhVZnD+big23tHg9wD+ne0M0EZkDQ/rRg4FEKe2G1u+uLwSWufGQ6OBDAc+y3/jZgmG
KsOjTuXvUqn4JZ4jpdYmLGNSnv0h/XXipNhRQ8A2PI2iPtXDvoOp0MHkiHtJZycZ8wDmxhKe4yt8
R5ZJ87wEhMM+87qlqTPwuz7tJYLOH1o5xKVqSbtGMDik0PyacTbdkiHBFpr8Fi9gZBbm9LS25hHk
vVSvsm44pwm16+90u3wLDuBK8XwkJcyVN2ManeZuZBXWP/FGHT8kQEtBTHix90jeeaRcLdoI8dBz
j7cDG4Jyhl2me7/ONoVhvk9k3Axh/0SPdtXcnti0coshTImkQy/vguz2uFcdHEI87gXCF6hJpTF8
s5q1O2iJLrn3cIwNS+T1DcNRbTLH3nKsajyOssGdfIZ/X09Sl4/fX+UuA/gEaak+6D0ORG2lOceU
u0UCg9FVa0B8FVUUG+rmqYK3jPAJzFQTE3iX7xp5paTcDIdte3ZfhHaeS/jNt6F9HWsjkerk6J78
uBtDA3GDOiRyza+d/VhSYvq0Ziw5hSjHNJ0/pFXleRkAA7UMW+4JCmCgR7/slh+LIpmEZiFPYvEC
XVuLDnbwe691eZZFF0gwJp0p3yezUIc5+nZ+2/UeiRFWrfihRrRndU4j6+f0cxFOwHcYMcjtCIHD
V97MUvkK8EbmpNaWgE2hF9Hen3Y1HoIQgzt9xB1l3JGmsQTp7uNtJ2WeeTYAL/Oa/fP/6L6SFdZh
oVHtKUkFdxJnq3UfYN6QcraOtqg9Vjr0IQ6vW7efOyv7RCbinrMmaieYXwndY4Z+uai6L7d9/jsX
rtxgczozpolq2brJukonxgB+TlXzirvTnVfFe7Cc4iJ1n7pu6MjlFWizRmDm7NxEuV30f9ZL5g9j
dtKQJBLGvdEVeULgZK4AAhS8dIRI5mi/g5+WufblkuJJDe06gqh96Hs7iNPLRCLWy66r8dUviqzD
Me5DVRHSS/kXLnldM2IVkXKWbFSOVx3hGqvtSq//FaJGMhb3zK3v4JMxq+QR6lX9vvA5RBDKwxIL
YzeyvmwTvd4Ea1j73WGyIKtTQw7dRwm1+4g5BfOYxLuR7nE9IeKyQ8dXobOugygMc04/1OGNjnG+
YlClfuPKvEU54M7hz0dWN9oS8thsoJV4Y15Qcukk1k3sRyFPhvfmQiQGe9q9v0vY6mcpkzgDttx9
Ijp6AJRieL9FjqGJVW3VIcAZh890D3e7pWkqkXT8FHf4un8s0lV1SUaWZORO/Nzr0PPDeso7k/+D
KrizVyU89lr2kxDTbboNV0WzUpVYAUkwDy5VVnam3FTN/EgZbqJs0DGE9783Izwkp8rUL5uRn2HE
v1ElbKi4faoE2veNySJPq3ESoCaJeNYT+nQIssUyIAyC3fNCedGlnnVYKN2M+FhxZGywOO1GiJiC
MTw/Z4GHraAizKmbk0gaDpw5DbuqPmE8EiJvjiXEA4lhH/7MAWrQNFXxihUz05N6LQW70TEfiNFC
qq5LkADO4TgKXifkZ4bVpslFDVgw9EiaZS+0UxOtFF+7/KesrwlYr2smo3DYYqsJmwbL2kG5e5jX
xnkbU8dXN88YdLLaXTwoX6c6VaMuUwTB0MTGUDhBkZU9CLlhN5S3fxNNkbADH0kp0C8OzYGLZIOp
9B9hGlKEPvYri1YTPrJ15xnThdAX8Xmia15Gi2ZXJ2cgWg7Jj19i33FQf0TSTFPooseFHX3dVHCj
sUGCSLgF7WXs29KPvYm1AKgGWMCDMz/ujnxbQO1rklu1on2Fi1ZAr06ixWd8g1Njka3Fgjvqobgf
geu6QezUcwokkdMcbBACggWpBsHkr2/jz720l63VwzB3gUoGE74AKxh9QZfzi9HmXwVM0GzXfEbr
BYnBcr1JpkhPikREFFYAvAGWNt8+kBL172O+wVVaYCL1Bsc1Pux/i5BQHYAB9W4gtAeuKcoK/F5S
7gDYVnpcYPf/1ec7VZBKktaQFwSWKTaadJE3cDf25BsLCSdY0VzjPThwuXhHeFesF63yrpHETHsc
xyRvkAKyudm4e2U7BFO8DX4mgnibvavZywBH2HPBqaNpVitxRryTUqXSQSOlplqaVfJ6/KK8j0IY
O6SI3dolJXnNIHtwwwdH3taBPG5fGREGcnKSN32pFe06Wq/6/Vii86hjtxqZvuxnSmghKbHVl034
F5Aqzx2IP4UUIXvNHLGe2/sWm4/UECIRpRG10vIgP0mEGnidMidZ8vomAS5uavSPKRKHyYq4Di0r
LuT9gR8oOhG6/QtsTPIT4omjDRrAHezBXsnZc8VH7yPhCPw1nSZaCCUhC9yHcrSr1r6wDmWzQUBI
ATHAzecK7g7VLmARfY2PHdVVYc76HwZQ2+8E14XWXrIkU54gjwF/cjKYi49s22PZxPi+PpRjrNTR
0ICbj19c+lzk1ypLI6r4TCUicXVJ6lpkrWHpCuQ/Oyu7UygmIjGy1vWH11IikNdmaP6v/BT2PmyY
qLh161c54ztUcamZCYO0pRIwIGHWg+eURowqI/il9fgj/ksO2G3hoWWKQ0C7ijUtkWB5j5O5708K
y23YV90LgSvkmm2xN9/2OmDWx49rqFrirHs1WGba88FIEsfEJINPFh0r/vO0LTEIH/H6h6FjGkBw
l1MMVKivJfP6xDxgR8Sp5Lg6N8UnahX5Ot03QeMxwcix/DDK0ifEshiihSxYX+Mpt37l5Y8sEd2o
Ep4KxnTvVyEGkPC44lVN9OtTcfcAAo63J3g/hlR2deUu9kTIGRvWTMhM2D0cR41DY3RGR+lXOsqD
gFDl/8V1J37w+Y0MNLSl0J2K29nQUl/m5oMwiLkKzNooUSWC2qUFk8UJlwKWRo0Cf/iF0dsONdL+
3m/q5MaGGQdbLQgHWWKshN6dqPZ5ceTS7tVJvEvQO5E7zY9ZMXpnR72jWirK4MrSC+jEekJ/UzRf
e+mD3blrlvQKOpULtgtWs/QP9dBupnpNnNCs3O4X8ALhmy2ORVCEjBKtVa3MY1lgcWU8tLP20blr
TMfANiRG6pXNqCaa4V7ewKyXuKDso0Gpsvjvw8Eiqne4Hp027Vm9JdWPEq+EGdMinoKT92sXD3EN
f41hfHb8WGOv6pHy2zYBIscHmP1mLQEhtjQ0pRx6BkcgIyzlYEQr9LBF1TRm/mMNZ/J1fqEjjtNN
OlDEczHfi/MGSgXmkxywcmNfzPvXo2b9Yv229N3U2++rqld2ajSViLrOwCFv7EFMx1X5/SDjDjXZ
uW76lkk1OzDGrC9qGZlaXkFj64gNW7uPz+srBwwVPaz+/owmnTv6D3Mj/H96JK2wQDM7nOafYyVu
lsGG2DQvUnoH/qfqqBRn3t+i62Zk4Kzl5FaT9G2sL31sniyapsqVrxLabYSuNIQ1ztvoiUrZ7k9v
MTtTRWrQ8UJ9e8VXK72EoG+Wg5k1s/2zGlE2KIJmGcHkhlzgWFSkUqxsNeORgMVUPSOKAJzQzXOG
Fg0SesKJBuL5ftvhMzHXr7dueIxK2jlYALO29miZh6oOvtThKYAF2UQb2XWul+O9sdZDYKze06sq
VYzzr5y+t6/DJVU5U89D6pPO3m8k6ffa3w9rnlaLIw1Fm1hdHz9zHvplVtMWWhXpL4rYU7NGNDcU
P/v9ejsS+9mIufiJcDelUZZHw3oGiXQcR3bqgHC7NlkAYKON6PlaA+Us+EHMcpclM0qX8ZIot4b2
A0iSYt6qX7MBZ5rcDgLV2KztIcAijWp4rK/kCulQCvx/AoHhhvUh28UuaZNRmw7pfQyx3csJxSez
ZxU27fxFcdbAnQocyl32dVaHZjpcarFu5VEj2rSl1wnddzEgiAkgXD9xeJQw2VK8Pa4FJM/mT1Bu
OxNKgjevauQOreCwk8iYnYqfAuAzYktkLG8dAcRqbS1E3m5o3K2nxoPlfoYtO1JGr8OUQMrgG3yW
8AbCvrY6ZYqZjDBwJk+vPJjq+evoVaRtcxbJ3YMSnbpJQJ03eqv47RY15dfvXcP/dMzwHOd3SZ3g
cjTU2mOFPEaoj/lGVvwmG9gFK+VWffBDGYnb3nPEf8GqhIeT4FBqPRo8ZhBG91ecHdDhfismx+qX
3bul/lPXt/4ieJtQhKg1wb9GcWqd0SFOGkQ5bNXvHgQgFSsrfmddMK444Xb+6E1yXL1WDplH7HT1
lyijJ57BiPipLiW+cw5m3yhVV7rDJ2MdkPbdLaLgnGH+k4JQ3XYZHdoWnIdQlKisc18DjudOkozj
Mn35hioHtiST7Su91EzvaMPjXc7Ky/bQAMLXiS1MV8r+xzN2skOoIKpytezs3VosV/yLTqx8S0cq
Zc+yOAwcd93tb2sPciebMYUNf8vv9f+8IKg/CJgLs9ChBN4DleQUalYTszFAun/QlXhNUQA0xtQt
hW3VWpRDJsAXR3Yt7WgpeOhszU9l7S90FYgiyJzed0uZ3QbhKpTU1425/+P04nd8Z3YBednFdaA8
o4PdvwW5mks3Ww/c4ssAisvt5HRpvaUtj36EpDweTAC6q+6nsJ/OTnS95dlnCv5vkHReSnk/hjYq
RzRvOsoV4VyegW0CCupY+1ZIt3buNQj63Ad6Dgzp8uwbt7T1Cos802KAXwH+lDams77AosOoBvZA
g/L6KdJPalDyRFNrbgWWyCcOWscsVmPltR8dmhawwn7cKo3npwxBSh/U8+CGCTCjlEi9URClqHLB
LZOhmiJ+vJMdDgdo7LZkrFdHmtw1swBK95xO4DYWRmfQcQ4oQuhhblI2iPHIIms8uCfQK3FnyUI5
dWH7W9yGZWd2TZOrrFVgpZ060ZBPqEXVuNMIm+vWdr3lZGjBVnMqB+lAMqqdJXUTNLOSZ69XcgWz
fUimuJb5N/Zr6OixJH0Gkp/+CkwfaxmbD3aMYD71ulG1rHYe6BeYJUSt/kYq3K1hbapp/bNDaDY3
IXvu5fzZFvc7tBLRB6UNiDeAqOwRGq/7WX6F7jHl0pW7TG13ppyF6PyVTbv2zDn24dY0nyNM1Olp
R7HSRiguR9RisxO9t6ST+Tg3w4FqE8/B6AK20bVWG2MuFgSJYrHsO6CrQK7dh8dXfIJxK3+O7yQG
LY0zTRs1v/EewDgloHLj9nDL1kM7RY4DaovztlLEgdG+kd3wiOazYpGR7lO93OoZq2kaQny5ZS4T
DfaScKp6m78d5jvMoWPN7DAxyRf0kNuGmh9aGwhg9hbH8xR3zRXDhmyyGUNqJVdcdqNeNPQJz1Bk
o7X/akajd0zGMf3slrkMTMju5oScjY4fDmghJtfn6LpquIAb+V35cmw/XaiO/5kMN6apx8s79E6e
y0L5fQIbMlUAx/hCKsarn9bXjJuOnLAwtIkUwvVOdstv646QgldiUEl3+UNWL9fpz0xWpMeoCGrD
q0YAkwQGWAKlU40nSZJomjR/VSNlg1je5QVzL9SClEtVERs44yaBCvPax3E6RGJ6V9UIrTA4TAnv
KFNDJyRlecoD3T60HfGl30LZ47A9QK8aATrezTmFw8gQhJToBxC+Jj5qXhuRnsboBFpMiEDw+7hk
wDm6PG2RLvJBuv0zojXTfJ8jDJUaPD3YOsKuslicjuPEob21F5tlr4MP347yMyzEfndEp1C3jIT+
9Y3ro70MBTJe8mDQBXdomqvqfQvh8pYQMYgKZj0wx4mOnFyYLlYQwLUlhQoDQE3MSO+ykcFZEOzy
zr6nT0bmrHPe2rmPTzYwnQyGNR4hG/9/5eHlVzPe2cZFSkBloAlRt7KA59IRPlHioJWKbcvUPtHT
ODWD/hEPK9qWWQKoSjdlsNWN8kEX7LtWsfmr9zcxpGWWRFxKGMS1+V4yZL9NqE+Kt5w2iJVJExnH
ObU64O8FDG9nKwwyl99gi3tUw/1YPM4Wj2NbtOuCLIP6Jg9l6TPX6B5MtHPMcDROfb2UhahBdVeE
DsPpEc5X64kzOOOkZfCGoV0RMqTFRSP+e2YszhM/VS0Gs2PTYc5El7hm/kCWJycxhjftiYYMArcP
L6WiKk+zZw1UZBCJqXl8i9D9n3PUbZg9rSqSwMEWPB0VZKEiDYDUzxm4uLlglb9BhWcEdn2OWcEU
a/jrhfkTfhcl2hWwHZBSIbaYVe6zYOxLrTXXWpllt38xL6swsxipImBbYFt8oRXTF1ruZNMsXtpQ
hT/L1nfznWETUmKfGwf3D2vMwvE/uW5elQpnquA33hbVvO5zY70AMnvrjhakSeJDbCa5qcYSYtu4
d3dYqNG+pzftwfmpndD5R+U1/VTbKPgWob4YRchSplHUeB+gzLnIR3+XtO5Ypk04/ySoBuTNTpPC
wA75wRGKePoeBVtZKJuDR2YmYA8PRwSMg2p0VF+B+aavaOMpwjpfqAVE6mu0ZsK+eOjqlKK4EiSF
yR6+IHFOKsB/X9i7m+hEiq6AWGF4ko1g8JJ3UbvdEqI1xgs+BwJcWqXj8Miig6l5t6ACNYvSQN84
7geE7LLX9ZHfryBsuybKQkeqHV7HAshd6D+IcwZiqo4Fsd3TOTgLwNrbMJcxu8hGnQdyP0s6k46R
XIAvGhX1HwtIgt3/SNLIagaWcXFmCH+NnM6hWB3feycHLeJp2sxq0+85/EeSnVM+k5RG1+rWGYZi
XCDh5ynZUcOY8EaVGkPAoVeXxEMGiFvXREE+OaBoBLILaidNRFnWcyOOmHD/o3hmzjBToTLLtYc9
v4OKUkqZ8RRTXPz93ga7B4gx6A1qf4m2ophvLUu/ZXdFiErbp+cEB4/jTDFN377UhkFHY1BIhLpN
eFbVfLdjyrGSvwwtG2Lf4xkMK1k5N50NK5WAmKz+ldJpnMige2yDA5MTUairM4hpUpIO2hmPaBH3
8yJRVAr5XB9jAWbGYG4o83hNj80xzRsGajstRVOePKKjUfhwj4IO6YKeF2kHX1p1DEeKFGRTx+OI
IXXOrYpAU6tSOGQBM+3Dice0vghaz+dwucgKIkzsVSHVCtC5HxqgkNWqi0FPtd6bK8LlVZopHz3N
nytq4eP5o4cgXVfWJzhpSvH/KtEOpgj1hN2vtNORKxFe6QYgauZsnfvv5H0gVHknRnGB46N77U04
tnfgWAZ1dl5S62BB85ch9RpDb/34TanxU4jt/2IoOEXUoaUU+m2xi19599202sQ8+8HJ/qUFSRim
ml8VZLIkxAsPcUYUBewHhfxJ7XWVaqkwd/AqBvkRQ7YHr8+NMC2zQGdIHBKHqxamDo3nGCYHBfqH
yDUMwDpzQBthT7l+DlitB0YxO1AeQwffb32YtOQ0QY8fINuN7D2JRrEDRfrUcdfEEKL68crNsMDR
KinsVXd98MvnUsnQBUKyiRSP3DcenR/iQAtA4dfIR6mN7vKQ8xnQDFVk5HTVtI5gypDkqmhuWTBo
ptNE5d5Ri0JIH6vVgtVj/Mz4bdcs4zJ831MBC0jkA6FdO1BJc8uOw78DoVUpkF0VdYzXLcrOsDEa
9mSCj0cxkZwFDW5ycuoX0RMpSt/1OnN6+q7kzc0En/uRafNVwMU3DIqQaF5r2gO6g5uwZVug8RTO
L92Ct/SOnENxEsRmQ3U86ISWeN9sp9yNW6c3M7KdY3mfBomZoT6LFuCCyppoBqRl2hRBVKTNre9V
kcegHVdFhMM9t1+POI+AtaAWc1UghEi/l1cEcnHpJNGAQZhb1ayBqIdp8LYuEnQX4CF2abUUJ7Hl
S7N1rG5Qzm/zlHH9RWRboXKJnTaSv/kJYruYCs7ku9+uJ5zZtEhb1n/mSePh5KgI7Y15zAUO5cby
GjNUrqz8nOfadCorHswu+nZ4sQPY6CxaKDpKz7x2uaSP6H0q8Xmi5eeN5dHZEw7ptaEQy34yf+FU
pamYTlry69Oh6/S/zalnFP8w9+A4kSWxQHKhv4sjAvGIc1eq/S2SxAHkGHP5SBoZWxIIvyBfdK8f
6Z6RM9HTY3hLiVGLd3EnQWEkLl7goCMYwcUPy7D1odk7kX9XoNYHUZ+M1rQKWO3HvEEGbpqW+c7n
58kD3F4iY5ckWP64V7Jdzdp1PY0XHr1W+60IhQsOsVHxIyR7WWVCR6mbbpfHCFHNtZSOiU4uZkCW
t+CtMVE2S/aPTnKnsIWuW1mgOdqiDQytTcYaksiRtL6eU1eFTvb5rsnJamCge8lJVJXEs0Lfaw4t
48FQyFZBRFWtX1KIlLXjpA2J4crwtCnFDpUJd2wcd9N+SU5QhBtIKx/GbWPqE0ZepFgo16QbVxUS
Cn3ehO0+G9mnRLcWhD00zsiNC6VB197XaD1rIc7R+bIHbQ8VAInXPvxGDgz873Wi0COGFFOxdZev
/A3K6nzwvdy4Vbp4ith1rV9Hzz3YH3BPsjNDh4yw8Fh1kK093mtlcOOGg8jYZUglPgQr1QKRXYAc
YZpI7Q06pazdJzL3oRMaQ1AHnDMwg7wDJT0Sdw+wo1MbTfBJ4sXcJ/ctPKmDWZfLu0Y+8InOHvBY
EQHyPnTjC3HQsnQ8B9otXAhL/zDkLwaMSSbZGojKqxWfbbvc8JKIAJkJGOyyugAHVH4NPZrPbL0V
PUGhfbbwU+jNJG46HtXNpfUuQPdbTbWGy2wc0nfd4XrwYXAmGqWBgk/tvIqnKZPFiYQ8vTjT5ZIn
KzGP4eMEAqgGOiZ7iqfEbqJGTkRcfmvdgqvDLhu4KR+e1IOvdkiSu7AyXX/7Jdyqt0Z8z3mK66N9
d738AJy3zraTUUx+oUGdkLRumteZshNUJZ4fnu/73rAmDseZyV8excPsk2Mi/2DNhG3v45j8p8Wb
UPiaLnxlKb7SiZD1hDuazLUh33dTGWAUO3RiF+vJUuwEeK3TMBDM7xeHIrdbbrP8UMKyIKm4aee4
CCjJQtCbmmOkVlLmvELy/Qa6HDkM89JoRQJ/PnFg3WjE/tfIslleqe1c5QF45O7O5+mhRrEYeF/O
voKxWQjHITb7CY0AuWsrY/b13jy8QfalJrHnUZT7P0qIcL9kGyi2ufBgHXDcbd4nPDslwuZyyMIP
XrB+PilAcuy6L4a9oTVJyWJVQT4u+lnNMtJIfD0Ic7n+/QlXRD/1s8A5TqhKlNIbGjVD9zYG1dfZ
JbPtd39z3TeC2tFLw76blTCG9zNH812on6ysLNe2nGpzxV1xR5fieFHx0gVPvIAJEstQ2lX+wSOe
xy/EeHuYqiKwQpOXlBlFXmihrXVxljxohm8XrfDV8xJ5f0jUzTSjUs4bLhQulSTMm5js4dy3MBoh
0aEp4aW6Wp2CEbru2xyGtyElHPGxGxIPI5CaBmCIfRoddwqaOZn+zwXmamoJkaZe19Qx11i98IGr
yh5/MrXLVHS/PM+u10jBauU2f9yrCQ4tTCE9MD/uK9fKdyTZvIxbRlGS5+dRwC2hooJtbcDd2oyI
KuDrlfro5RUsY2Yv3SH9jm+yg3tLCA3MOV8o9mMZTyRwXjIRtvh9H30A4hXhSEkyMuKOr7CnIoCg
1DXK3i8CDHR4lt50Qf/ok1oezJ9cAKCwfYpjXG8iwV+XuFYjen9JutaoCLMCJjvKPy5IV5Xp8H+J
0xoyLNd1qI70PiFQOZTRp8akNKZCEivlbCzqap16oVDQjRQzqm3psSszY0kuXvu7hsvI57F8wemY
8YqDExSBzvMxUWOqCZNv64Ej0b92FManK1VtA88cEce+VSfWWMl24wjuiaapFAtspbsGX1R+ZXnw
nBbk25dT5ZeAFiAfMdjsebOHsZqFASmZP32aY4TPNRGVM5rkgG6Dw15++G87dfSQthel5CO1UK8i
msuyLYRFn8sxcqZVuNQ6vSOYs04Btn2ZdHcRk4HeTO8VPuPz0MRYN6hTyUwAH920bEAANH5O7bca
VPIUHuOwUcRZuTXSCudTSEfRRB+IXd2EERhGkQHdwoBIzrB23mZUY7OoMVYoKcvxAvjsye9dxywS
QDJh/oqXBuisiKyM+sQZKchVSfSrNfLa8W161qfBYTRGR3iTsF3UEXx4/iCkZNvGTsJA/qOdQe1I
A6SR7P9iXdSf3wtP5YKFWNJZj7xXIYUft0VbDwKhTlX5bBzyWclH9SBa77F7EUQ9aHi9KCEVovX9
/HatcYPVc1HyCKlMx+DRM92YhO2UbbSctJag52FLxGXN3p3zqJvXRMc0ovnWJXbm6iZyGc7F2nRc
KUD3iwxzCajd8T7+erQlveKf5ZRMzH7e1gVcI3+0SqPV4rsanAqFLWL/Fz7rkk9CMygvTlk7Zx9V
eNm2jQ6u94vzbHKR41nLd5a7x6q59vtg34lH1mUYklLCyiVsao4rL2J8LiTml+HH1sWqeLkYYk+a
Vjmt5v48Gw80Lx9FOd5/dmLJ/lvamC926+6lpeJxgtpYvkvC9Y/MIAPuY7RXS+oiJ3APxQeBgHLL
CKKGSgd/y/DFDPLCrwmDIA85pNhRCbW+dCUwCpaFbr4ldlUmDd/W3YrMSv0tk74cVyD5FFuP8IIP
QL6fdvSfjzNwh9k5gGQeuJG6HqqR9nUVpjJBXMr8VNV1KzjOqLj1eWKKCneoBIaLC9Aae+laFwVo
+OBHKbMynACxM6TYOrrzb8UGPvIeQGoDBlVFQIvjVHh+ea7d5T4P4CdKn5/+Ljs83wyEZpQSicvo
UEOoE5Pb6OvTy9A+53s0W37BXL31VqqoGl74Bkis6szzxv8drIi2H7kBPmW3FalFOJ0n5VFk4kHi
cVZTMV8Qg8fTft7bGOsFQUQwEG/TuPCPv+gPVy82VZn2Dl5ItiimIbZp9vb2Ef79gV+wMO+q9BUq
f4tc+U+Bu8GB0yAekMEum+V/4RIHz6Uuon64rac5epaA4y/D9rNfSsHzD0/nZMESGsRzyFrP02Cw
fOrFGb6CK++Ba6czwfAMlMO23bays7FgCVnOzdRb4ASFYsl9VhB4esOukIyn5LSEiiD8mT0jyror
US5C6s2xD9gbdzvNr7VaLa2c33Q9X2kKsk6aDU0PavfZdsQMCTxAdQ5DKR48zU7ByQP89tO7YwWx
fW8hRL8fSkEWHq00t448Yn0cMHLxjFyyjMBuGvHtXyd3YBPjNzzWl0JFLV1uyvZ8D4YgfIHirIkF
0mE36PxNKabTOoBhfBTjeo6OmEJbO/Tikwz/KdISWRU3n53AZsUaUv3+XfCfUPxL52NC4aW2BIhU
055bd1n9bHCfGgNUZRc4+dIEyfvwcQcoDxsDhBSY1OKJj1rvvxwjlrQwSEltoCTTd6SXfBqD3JFo
ZlKCwqxJVOUrSVCRfqC62zbG5EV5hDDyBENGbqrod1DHZ9kdtf9dQzxxh4s3AM4h9f5PRhVVhu6Q
3JnyY3fi71gvMXKzUAdiXN+CMXQHgkzF0ej6gTT4N90CttZ7bm7OxkIYS01Wvbjo5Q0AJjecmx9b
TrivP8jplori9DQ0N/KXJ6d1ppIJoJ0YgiJBFrnz8JkVxaHr698u3a1Mi1pxPlh7+ZyUqbqg6M+u
jqrayp0h4X/v/08jTxE6i2DOkbDwCX0TiLXBfHo99iv1fu3rku5Gs3FdIdkziieKG7nYF5E/vdbO
KWof9eaZN2HyBriJQu6ZdPJxhYn6YRypk+kdQyMoku2FKkGQXkC8S1R3pQDOD8utUjh8oCXNSLTc
I7kvSXRJ1Qcsn1IjOYQVLLM3sJH7HrRGq2CTvcr4ftCY+DgpdXSzfTDudUNmuL1hmsL41Yho9Qnv
I/phJfrdjpdbaT/fQhchunHxe8FzkZqsVGVZMBH8Dl07UM0bmaoXM9IlHhYadqDjvXcYpLbwrb0j
kSrG068nZVwpSaUXsJ1wZ/XUltdWvfCFTk+UopQXqWdFSlUpGJrfHXVtW+QMSUbk9ORyf9Va9x3u
o0lZApI1VSmd+tPj77COpPXmgUH0DrNG9O8TaRCTlz6+VHgxZdMrUZ2DGw7u3oX+eOYXKlck5M6F
6SZy7Xa6GwvttKMDBruejfZIkglPpJV4GV7qdt72b/2fDJOCt3cI3o3Qblp7be2grVKyztjutSzK
smGEr8iciTU5AP3d7Y4Rkoe4gAMs/tn3iCmtAk2sRTlgeRkSzpYHBmNaQCNUchuHpXT3k9M5RQnn
vYh8uGdgiMmD9pNJWYL49XKbMuxZMiGhtZFd0MQdSJJ0Eeon80AoYlcoZmmEzXCLuY4aLLPMtZnZ
DhbfFYML0eBQP6USXNSv6kqaOUq0wXUjmvx/slLC0hSELsnExDHo4plkeH5B7t7WSs67sF1usD5v
FAe8XuLKm10RuD0/GAja4j5CEfLtOGzUroa+OdXUOeCh0O1gPoFLzrKE8EYqY+zTWzyZhoiAGBBF
KFNet8CQtXOqFF/qJ8AFZ+quWKWCUR8YFhF4ezoQ5Ab4tReQ0HzIpWfw8uyCBLzgLfaor2YocdW7
hInIlnDe5yHAeTMGxd0aSfEbafbDhvunYAvDifk+rz2+xFA7myzVg1dCtKKXnLDhBtbrzSbiqiSG
FljxRjcacN1aB4E+l7efcNCzDTF20CizmfaMBqvH4jgCWf5Y6p9muadKZCzuQmXUWVpjrVDxf577
WvTllwOTve76mf1XPJ6lP71JwfsWjJDvAgJPDiu/EXmn3NvpFk6cdTPg3NY/Guu4e0VdGckq8IIS
84fPE9HfYXtNAFlejKiGTJ7CUcOKxxHaWDTMOe38lvlCTD2sjrNJMAJCvrg0/hNSC4KfMExhmH8S
pfF3IK3lV6eGC5xlKBJ6fsnXwulDpNBzAPzBBE00sefJr+qy1syn4UkkRm7CGjqIaabxF0h1o9yt
jGsS9m2ZTLXdTrr/f+sSadS0x+XNaWGS5sVm6yxNeeAGpIhacwyOHjbCwejqy5ZfGjppeaGBToKX
EFe/Nh6XTLbHIccvITpBTAjQiSNAvSog5S2SqE2QfrxN0gCLGnLbI5BSeNYK7Yl9KFY4sMh0sDug
6h7FWImTX5r32JKH8aazEq+myMKdLdh+6u4wD9UgOkYzWiB6VjLzNvmjmd3p5teZU0lBgu3gqKJx
lbiuTlzIDHrHwXvVPFdAw6S0jmpZkSC4LpMA3Q+lj5+UvfSShuKQJArtiNRZi985F295GIwaadmL
yzqUOX4qqnuRtpvt5rkP0+Pa4MG8fQlNAnpfnOtNDs4xQiKmud27+Li5B5iCMFPbiNr3FqzSTQys
I/NKpHddTtW5NIDnKn5Ns47b0wraRI5ITMenDdM0ILin00/9h7NF7LF6v2ndkX8fHkaZaSsgk6o2
JRToUxDjRptXr24mfPiPi1OV01q0KJO6qmR5oBHCr6D2/2FiC0gKEieJp2OtXbM4g5eqDgLL4oXv
cuJjW8Ieabj1SgLJqgrmrO4vI4dKBVbaYNbvTT5B+88c+B4jMdt0ScwRZYojSkgHUmc83OQzyA4k
ZUSvLf/P5/yz0C/F6QPIBpf3rE4u16FarrVTQXwUzUBx0st5iR+2RlWQ8goKeJDUP3rxWurf0jsU
i9eZG4Tf/hocqqKFxYfYwgiM7PuHvVOxQRGDqolIj8P5sLXNL5Q0xdeZOu+tuRLqf27oNPrQC65m
QAEfqtltFmf2alwQ9udDVE/7C4yh7yxMw3+aUuHgPU5dvOZq1FrdldJEf39AgMNAlCHl74dXFbf1
/bPvc2k61t8cN0ADBOHBrDyiOuocIK3AHOG/hOPQWEOROsf6nCD03lxK26UopWd90aow1r5yQA8v
fJuARpqAW6VcXDDZVI6XkbunGwTiORTsv1YbKp+h5Hec/DMvkgjAj0onL1S8G+YzpNr+HcsI0Z0d
M6WlpWZyklHxm7GoZx3MlFbVpdU8DXRMrVIhkUHHrVApxKvdkOOkIw6GBKdu7Gav/Nopgr3Izzq0
Z9lJ6AmgB/uPnpFEs2Hv6shzRy1HCxuBd35KwDzIlKKs/xtvhQDwo6b+LvGitJFPmBapi1Ml2DvB
GQCnKrtDKbUx+KL45Yjz3AOkrEay/xY4+yFkPA9G9s/Jhh08QZrOsybgu3L0UjVlGt3ZDE3Hhk4m
fZQlrAo02NzZFSU1uwfO9f2q4FRfmJb5KSuIfT9EuX5eqweVyrSYfs1v/4joRPqPl8cBTyZIOfZN
aX6hByzKAa5iw4eV5sqnnRvYqk1SGoZxzk5xnkUCn37I0ciT426W5Exsxm1J7aBx38nKm5FfdJkM
rKUtvY8OIzpWMDTKwJgNzzX+V2kiis/+t/PYWxfDqmSNxTeN8kG4XPu7Cvnpnd+3yHOLlfJRqMVM
nZBu0TZzi/63OQlrOFLUxwbIC9LpMJdhYhmsjvsAq10zG1jUYbyQkT/uTeRiDPJxRw4lg3aMqWU3
NUnunxY1qUvr3HED0Cs0MFr2j0NkWR+k0vi/mW2rgcrhbq4Oc3o0e7RN05a7QM2VsfGR9ayopg84
iOnO2x4eulTJIcspQMNQspXy1hGV8NWmlILBE4dJrqlDMkhrIPvL0Ix7k1DSZBsA+k0JyTgcdPzr
DE9ilrgXTh3qs5z8mg01PcZtPgBbWZmJf6sYaKinbCd85jRsw9YWOmkoCzAs27gx0B3h98IayDo4
DNcwCai9B4Zymnu4Cdl3MJbRFcc6Q4+p/TscEY0DZXqsdHaAzbEHhAvAYuUQ6ODr4E8HuPvMiSKT
kko4wNcfy08BU9acO5z0R4g5F5QVcZ0rt8KLq0eSECnbH7oFJOK0HbelJKAx3f1aZgIhJ9WrM36i
lqhHTbdc0jOGL1itwDPMp+3J7yVKzY8nbr+RYX+IVL8zgWzMe1LShYkyIt+DA10VpPfBDCSEGAIK
EFgBZTPxNQjt/0GU3f/bbONznIQgYj2qF3TkjRdDMWHGshaTCFHkvYRvQj7ZwK7Hztw+Mtgb8j4P
FskljxWg3USShSFLXdTfJ7IPybaFnWcm3Bgzo2DneDEgVTvYVi/C678PFBdl8VQ1Ke2Or9fFxhsl
lCMK2jMKeD0b0iLsUP8KPxCS5GZLOLAbJ/LEe/DNKGq0TWcpvdtOt2NvPVAX3qwoIhmAu4g1oG11
DLtllBJ7vxf5HONATqffJznHYV/4pLAj29xUjGSmOn3ni3GjzC1jKRSRYowr34nBxt2WuecJQDwj
5fMD9pyStGmBsnQc2+8TaRAFxawPYWFg1+JNxc4wQV/E/PuD6PIIA5ib44IVjYZ3f2LHKWRBZqhi
i2+ZnMd4RpZV6QNuFypCZy/TeI3wBjPzz4YTKP6m7Twa2+sLL6qF5EbgMGxBfnRSOjy5zhwHI2ne
Owv0eX9AOBswkX0yqfKPtND9ro0TZHg3CQ9rrmnqw0cdIX8m3N7umk3kAV3UnmNTCj3GPGbBgz3l
jUoFZdD7VWt/Bv+X7geVr4RfstReR7anGdMu9FupC9P8Ik3w8N9HI7kuhEeGlynRIpI+krRRdCSH
3UijKiXYeeX72osax3dbhO3fUlWVVLBsf04zUJ3ddjJqN1Di8BSHog1Rq4Z3r1H4cHRCwI+hoB+p
OrUKkqUN/S/4FqkeP3EN3BGHCEajNo9iymVbM+VTnA9zFKxwgubWGSq8lNuegCH+ZZmGrIeGQBbd
IHRR4a7ESAz8fi5wNbp4JHlzGy+BlXto7uycNtXfixZYSfF1I8uXbZnf5iFNl6W+nbPNpeSUDAzg
/NqDUfpppQVB9qdMBdWhzt6axeerjLGr1umFg+1c44nVaGKRGjqzvyyY2s8uiwlE2vV477FcfknZ
tGY0VEtrlKonUE7dRlkcph/BdB6PpEIf+ipEjR91BvRv8lx2JBP1jaGie3xx7TEUOvFLsciWR3HS
2UlRkRyV8Y32tslM2O9TDDHi5zDc+OMPicXjb0lTFMMgrG36N1uhGFFM/OVKVZ0QI652xoyTrkxP
TtVCfojU2Kqhf84Q1HQ0CaOtJd58FbbL2US/GBbcHpqHJSJNtPwDJUOWUSAVH7L7lBmx1p0WEvNn
0CBcOTdq9x4S1Nj90C0GP7K1FM9PObnCpbhhzIMfqzUipkXtBYDKOx4UMX6c54nR/NjQZAgbvDfK
/828Aa+RXqpyp17FZ2Z73Uttqjbizu3nz5pKdvCuIipPPt/faGOTpUCEIJSusOQp/iyTtr+JXxzH
f9sMwUX5mO9nPLcA3zo5GHjtaOgsTke4xTqID6eFK6kEWipQZFc7ai83+eDC8HpNaWTBKPK1rFhk
69m3YjR1VtdaXLkw3HgokVk8e80KEMcPTuhziauAMKmlIYOS2PZGpcXt1ZxUwQ+1oR90T4AlydVA
KtS728A5H3qizN0iHMS5lDkNi+PMd75vwIGytZFHdwh3p5OGO8jZXOdq/rA/EGbDdoa/Yb9Uaf0+
kpAMdrud1yP9H84+fNl3i0kXJ9TwNMG8i2AlR3VxXdgmEJGBxf0toD/z5LioBbNAYNUt/oNrB4zD
yo8uHmTDwLHxO7VMimLjElAkszhwL0JwHprpKaSZ9ToDrlWSBh0S/wkvCJZjnvlxXRf+o9cIp0Fq
9m1o/D8kahKwzpI1okncvJRMTVSTejn/Y8sgLRry9XTk5yPBG5rC7J7DIWykOsTexYpVHkGBrTAA
r2G/DOwDn/Zl6cVMi0D5Qb+4yo3rfBnMWKrRK8BIj6wwzae042P5O92xTTAyxLV0+1H6QxNjpjoW
OO6HtiFFei/9m4VBVIJ31hG+Bio+YaUv7bMP2jL53Ie+pCdT6ErLJT4x9+/ZWLeq0U6Zn5vpCe+R
E/8xTjLxNEbpi8A7dau4pX1iDPb76/gppDUvmZA/A10hJ49wQYI5hU/dK2ui3F7lieCdxLXmp9XN
l4FMMoy0OI02f0sbmG4ack3f+hCiOfXaI1MBNnuBIqbvvyI7Ay91Hk2/ax+ukooClFiGFAHn9CxB
35MeKs91remmNKjyMRfJcipiyKwdvLV/Mx0ieDPjNu74TsMmMmUSTXJ3T91yJLYv8+1rYcABwBDB
yD6O2InlXe23OFSEzdatFulBrxMGLpDEjWGPVpj7fwl5kOLTWscTYdCtb4v6W1G2knLVIOXmg+jD
5g4Y//ThGsC/lekfbvmRxBp5Ih3HS0F93p3WUaoIDECrHJGQdYVg/xuKQnceVFFrux1GKZXsf1Cg
bJ27HoWZAbg1QWFJMgw7OogarbXfUncM2zxEnXzKCMimk1LqvQ51qVC9yCHN9mOf0kPZJULuqQKf
FhdUcnJx0msLTAZIaWsKh5NSAfJ3wqulR5I+84nc6VEZO/oOWV4VPvU1c01VjZwqIjsdFQN+28s9
BAkr7PHzJc1xb9CmARq8hFe7hYbDCziGlDJrWIfQ9b7mJR6I7nV3vL+6j87K4Aza53zeHhKzaHO7
saLNciErbaATKRCV80LpVG+KwESwb6cxXKwE8PD9PHW8Rb3RKPPoq8K7frkm+aH0M8Cy6bykVRFH
KD+wdzlYWVpiAI1EnKYK0Nxe6RpvT9KApADeVQuPaahvOnRb/8G+o9+LWHJPYRawE6jmEbwntayz
sTYjkyQCKqwTd4jqbC68a+S8akC2Lc3ZRgnI6ZePMjcnlMQb8WrX2abarNJn8eV3iU+L9krdt7SE
E9LmsA7ZPNZnGzBBpUYecyzOvHfBPlZMqVp15yfM8tBnAD5Z970kRvD3+pFo0RbIm5e08fWX4em/
k2dBt3WO1RCW3HH34hhFZJgWa/rnS6GzaBHAdYv5vECnT9u26+uU0KUiyHhZSPKn5RYBSeIoZGxG
DhZXwKS79AVWOdI7NC0K/6hRzvFiJgBxN2sVKYkxgydEj0SbGFiZ0zXsM3mwLuda2IRSq6p5m1IC
YHNIeXlHINkjpQH7N3qCgFOacO2aZOsMnlFXHfZoD/M2FYDUh6dLbwqVf6/D1aTr/UZSIXroNJKN
GENZ5PdF9Qvo5kJ6RkYZkou6z9KO+6hnf533uoxl0l9ftcaehZogkTUoMvjwtvcfrhpveFFmnIe6
tSrQBVf64lPaE425UGzwrXHcVvr23MRbRYGidKoxPIlB25IVJRan9KF3tYDdAzgXNR+j5o9Ju9Wv
hyl/1rEVfjbtkc0fpq5nN49HzMDsB7iNs5LiBrN20lwxKwSUcXRUqLSyPO3tQxMFeWH9aJudNsis
Ap4nn6mx98GIu5oPl3ITuqMO7BGioywbxZTdoZovkMxA4oeWHDyYWxPOpnuRcXvedCF0aFL0ErA0
a3/ox+SvDDVKNuZGXnXobD2Z1d/emcraOXzoq07IGu5S8T8NQeyr8x1VMkd2H9tbprs6ID4XilMx
+d5iGW7pW6HQiRwUzHzBtc+rSZQRze2kAy4WacrpBjdmEWiAStCNVqiqKumxHDslTJaeS+beM/1O
1zY5xPgcEAuQGWnxLB+qgD4dOYbHz9+5HUqzGrOmdqZsvE7rfws8yp64j82/3Qxc9QN/t71HtmZl
Utw/jlQYxPUBScYZM80PqZhCMT1tHtNTt7xO0N/U2U1QCE0+UBSXwx9OgA2Bgw5Q84qVHs9zZYDs
wjimbnQ+YmdPc/BCo1LjEoUsraqtsSBwdgCqYthpPfusI84MrWoCEU+bFSoVrev11/wLC1NN1cpb
VEE8QAhlN3mwej1FM3FP1E1+drBmaxhA2IrB+zQHJuQ8wcjj0cn6ZcROYghI2vtdhIf6472o0ier
zYErJczh41+d8DwoVBhP60/hU4UkB6Nfgaih5qq3uSV68yuX216F5vSXse24cAEOP++PR6necYTq
f1l3btIMNwBLzdiL9muIfnVoadUdMdRub6E45TOeuECtgr+4Mi8rO4oTqN069pvkS7oSOCDf/S0A
o5xVn1r2hCwE7Q3MKEIWi3SJSYvalYTIqvkZ6Ngdj5YG+dwMdQ4J5xgG5/7x1iLRJPqq5G/wf5FN
Iox0JZq2veTww+Zaq2zyq27r4kfRQt0d8m+shQXnr5JYntsB/Cy5zAOivSQBhwRDmkNQTa5j1LIo
6MkaW1WC3irb8a5w1ELzutIbYW2n9LnxL1Vwd/kVPEqsqYAnfu8EZtLQCsUTShHHcDcUaV3BJ/ol
GD/9+ZEwYEE2DjUl8xX8mMmRbreexxgs97hDbbz4PHmy0/kGgTnaZTK7KtyvKAAs00r85zLLenr/
rxIdNSBTFHSw5uYsd0qqZ88vYHb+dryC6PxczPOb0caIg/g6WUJFBXx5QAYl30PI9kY8OBO3Ce54
3LX58iWGIfhI8JoaGOGF83nnBuee2KGytze2WGHqR2j7fhXy5bpAiDtJG+eWYUjRTEgrn3iBUFES
cSuT60vALKOwLIX15KwABcUyOdxenRCdQ47cNIMRJKvLLNofd17DBdCG2DN7XILSLaj+dSqMQCTZ
jRTJCKDxKce25StwdG22t0Cq6sqjrqcYLrDbNjOcUHFk7oBUEDWHasAKsXNOgpfoCMfX1shWNiwN
dPbyAL2De+4hPalkdVhh/cBxvrNZ1roRCuplVn/QrbYgwaR0Q8UC21LYAmIJI5tcYvL90uUYNuBo
Smm/MaF5W4fLH3HKBKzOsWZIkOxGX8gqLMO78dQuwg8XGlIbWryyBJoChfiJqDWarzcn3zNfRK1f
XAu2zmkKt3jJJuslCilI47JSQGfnOoe6/0q9aSut49BCcxtN2uZoh+ILmFmOtkXID/cyTJd/ttlY
JoS8idxqEwcQ3f6Yrqacz8RviuE86LsZbgxryc1um10C7x95yO2HjO2mMZ/QDwxVSO+TlI4n6K4P
GW7MVotmvoWLd5VFIUqqaF1dFCiNUrM0TQgWh1r3tCVaTkL2BrPIVXV5RNDj+miHY8poiEMXcs5a
hrie3QnNkQWd5OH3JKsOiSjBGMxc2kTc5/TF8XI3+XpBHwOPCfYQITVFtxkFjvlKe4pF+Jw6dbrB
n5H5GoOWu1O+d4XjfGcC4zF0zXKnULrXhM4iqUHtlFWkr8TTif09jWYLKw5GXtEfjKag2YbF0L4V
aoV0dIjMeZKK/GMgC3MTwbU3UuKur1pvF9rzcl7PU3xz9HiXnBxcMhh/l/LeQ7HR0KPoFlZNNqUO
DlFCM6tQSGj1gWNyuybt2Ei9hh5QtFM2D7YbvSL3+RHrv20LAVuaTTSwdk+uydAo8O9cGDSv2Q3c
AuBsKOR75i+CRmH/61xtYZtZg3ReHczNuI+52Bel7bphq2+WP58l0c7AvDDt9dMpoyP/Rl5Sq942
hdnMiRFSlU6+2KAthcjyRQGhJM3LfyCYR0gDHHa0NQQ9QnP8dDYwFd5uhhaIX87dFiNQd2RejaLQ
40yaRMT38R/G6D1kHZIu4mk9eyI/2fGAxuvIq3mZW//vHo0nrc1eZRIOBxitFG+IYrXP7Efzthvv
h8ueRm/ontiJlVun7w954dqDSH0V1u3C5by94ZhTAcMbI/FKbB7W48eKyWhSBCEBKjx2pzA6wjLv
zX3AyDblcfIFncufAcfdE/ijpJ45t/pSj5NXmzNpJoAzsXgVpDyi3fbAp0lLt9IHN612P1adwV3p
8LQoCzxfKiNIRs0voJn7aEnJACWIxiToVG/eOvuHdZbuCD8CCGe+Csr4g+gUCN36NdlSa/zNrvk/
VS0drtCOl7lIjylwx1TQMTX7je20mMILvNvzwDWgJTdv1u7HG9mytGjNACptxlWvXp5Os1LOmKA8
BfnCr48RWUGFMaqHhHynyoN1Ufg824dATGYc4irpVsl7pIJujNTT67frYUxmfutxThb9E2mC88Yv
TEIFj/gKjIoULguRmFQGHJF10ky+/JHuO7xLE/0+kostlrw2zdYZWdI/m3IoKsVdmyQC6x2mHzGq
MTDhfeFEFL/y1GAzTv8doyLojkQdOMZM93NdMyFKr9n5LPuJXB+CKN/C6eu0BQhbBzvSy6HJtIko
LjBneCz6S/g8sh7GQ9PehBpMpXkGf6YnJ6KOSHCM19lwUrmZuRpmIgSOxQW1jLCLqNy3YH7LVeRA
TYTgrMGQPu0i68RgIu/ho7xNju8/2Cph+WrHpuBGc2EKTkW2ztdhaFGkQUAMle76n3cuUqCe6Onb
VDymOmiinkE15bVwedYnnu02iGlsin9w7EYk6wMCr9HfFrphd1viL3G162yr3EfBPp/ZIJosuxuc
aUXHGImVGCe9kb0DD4fcI+0ZCFH8/lAaYSJomvax+2WVATeoV34u+Dkp/jRKp/aMEkJE+wkRzzxq
NZuRIZLxCPD4r+7coS/taFQvdlPAcwfqhc89qYfhG3scsDXHC2EabeXCqLDXTmwemIFjJzYqZavX
kbqnA8TIbJlRhrpsXgMNoADLYiNq4zVqG2aKuQ3/MnQ0Q1ISws/VCs6v+P+6F6fMU+hPMXFQku2i
ni7m1npqfBVqCiqrRrz3nLoCdaFoO1rbVrPq7rD7/oSKGDBRX9MoyUOdoxtNvVqg/paGA7ZfQhqq
exA8gHrete2esxyvjfpdgzvhvaCN4Dk6yhYFYegbz5Pg9FXq+wB1Pjff0LD1/wAFXrVWJMLvwCB5
nuh8IQnVMnP4N5hSUABeDmF0KwTD0jJeGzchvdnTxJchWIw8AqIblgWbaUTxRqWy1+aBCV9uwbJx
M9Bn58Hq5+3vN1I11T43Nd72ISPXx3lKY/Hw+DOWRCZ4iuOXmH+VyvqNiP/WTYPLYdlz9UATmdjf
iJ04BSC2nP0u1eOTe1cZ90J1FsFzw+f6APksjY8hPirc6KE21gQlFUOwgt4IHhCZ7qswhnYOLoqw
mk2yChDvQ+BlxNngeUUQYhIsSGyax7+Y6ZGRqRuaPM5vnfmlGxBi62ms1+KOgFLjfnSD9YrsxAGQ
dg4W8FJbsWsdnCzmMcMS5v7euFDEGEE/ZcsPkWfwLwCUgwPBtS6m+vr+07VydRV/RBRFFcWtMViX
pMvZgJv9BAFf4JstbXgjXXTk0ZIWOmG3bHynoTv3jknqbnweJDtzflzUdWbQUiPq3YvsISZwUtgl
toD2Q6UL6X07kG04CNU9wgkp2UWZ2A1dV+qD7zQFj3945hxc/nSW/xlcxfz5x+FxaMBbdB235q0g
zQaMbBsdEWymSt7Px+2/Lw3L4cu7IIH8fXF/8gkxpR4/ST52w7F9nC5sqRmb7XRhAky6n6GmznFD
lrwpJwXtnwZzKNkFekPWdBo0Vx4yKjxbAlQEncC0/75cHl85RtMJNXer2kL5M9LQWtz3n5cApQT3
4bucQSGBAB+36aque4IvxcRhq0nJQ8t3PMDaZdFsMEY1avZR4kptVTwjrIYA36rNC1v6UmuhM63v
EEkW7fLMtuDb/A2ivHsg7D64NYCvb9CIbYVjr7SYE5L0OHx5zb+lyVgST157rSyu9d/Ci3oQl4kW
T0mJGMegHLEaEWpfKBYXT4z9KffWIyBXMT4Gq4PCAyz6R9wBk1lVeLCcMo2r+vSHp0k//PW5f1gD
LDKasWqD1+3/PJbYOclHZ+9dDFhcyJmgN4RVDWE3wNgG8Ck7tRSf/A7xgvFTk/JP+j0l1vkVHb78
Ast4UeFwZrRh+do6DVbmDyzmty4w5yOnPyPUfRmVCkpN2hXkoWOBDmIEPjZr8kRi03NwwIg5qGDg
fCdVxeOm26c6I4b2Z3f0FynFsGzmvwHeHeE1Fd2SN7HKU90efZGSdz+U+e1qqAHB0bcHxKl2tkOb
nKSp8c7vsR+CXZgsUF8RU2ASWkQZC+PVlf+dNxezqh+7odpOjmBoizCiqnDlyrDXBDXqYXHMaFP7
A4nl71uEbENVMyeYOl8wJCfzJRmXjJcKOf/QXoS65Og5L/Vs1EfB6fD6GDaSe+cW8t5lmhcieM3G
hNJQs4e4TAvayS7CjkLLR/Cw/SoyDoWXx1oT3vFZY7CTGNSDSWMu556AbJvZJbjMKGF2qOK5k61w
M9QNX74xI1ZTVYJTip7ZoqzAdZpd4WUlynYsJTpcHfjAEZjnkeQ+QhzLzPxdtYXFxNnceLrf1cUU
qLMA9a3C2Cyy0v5i0RvVJpz4a216bzbdjm9CEkjkXnuahp18VNzeMGf6JlZ8H2Lsqp7zi34LhtLL
w4qOMiuMM8ixMVIajnUv0h9jWBZYB0/sZUnvFMF9jR8a7tJ+rvmTaCrn0yP3HeYysAd94cOM7z7O
JbyFPmYnXH4gjt0ZEn6FKKcEXOkl9c+m+grVMF59M6p5mqtujUit6WxdLBCUE512NQcziLWqObT1
tnocTFB9Y5SCGojT1FA6RMXRIzvVOg1eKFsJNCInx+93GK4WLv3JzMSavWUn8IiK3lOGrwMnQExR
IKZoWrmGshXJr4YSlo7n/WjU/19T4mqXL1UxakgqpwDZ0sUvDIc9nQc5a9/zqiDCjZuJpc92RZCk
IbaspwNL8Ab4alEljiXF+vaAX55Lttzebu2CIlPlqBxFHCEuNUa2Jtg7L7HTwrQenzc8ur2R40hx
bJMuONtxrsTAoDDSTM0HHODuzgX4IJpkEhQ8SW17ZfQMazI+ysrhLn0QYPvFLCeDGr/EqCwwz/OR
wXj6t6Qg17NPRCZIutC8cQJXJomYUftZ7pRcFuQAfgsNRVJXnUejzbWG15uJpyU22Abu7eiVVmbF
ZmUiFLgnIqP8ec9DpQ8e3uKn57ZHr402k+ZcriGUsMRWHfE9/vL5lZGj8WQLt3LK0PuVHFYeBNmo
l6p2HgMEzTUDaGbkJ7egmux28mjJwx0EEOKLQ9vzUUl9qITZ6rlEykOywRYaqZ7fCKqEQ1HXaxJM
CBDwAz2i0QA1naz6xdQf6FuQANl52itxv+SBVH214yQO1DMzMF1y4jVIUHuIqZBR8Pk2NtAATwDG
PR840RoyuMAq41034CWfgf+8EljLruNGbFI6J5B3ILWAOhH3/RXKe7IcdcIZMPUAf2pntDIFRQYr
WgdhnZPFwaGGNS2/F9atgUxdxj05NGBiRwFm7nhi4IM1YJaHVsfTKx41V8NlEnBGClfDXUmYVrcF
Q8eOI+jvxJZ9HEgDHCw1z+YEJonjMvxdPGGobbHDe9+ZgJvNvZCyc8tSabAoHul3YesjpdwZbZ1V
KNksK+ilyOWEV0qIFi6lz4JrJL6Oz1oZ3DF9W20TpJSEV5DROVG4Rz/oQ6u4r3wSbP7m+SCWdH6W
udEtQpt8KjLPUkBsSXowy3+2d9wtZBlhIylCajhZJqrvpvzHivY79zxyYpJdvCfcM6AsyOhTAAkW
VPlB40EAjMwSyatdLbAXO46XlxhseA5ELe/VaMIaFkEQcljmu4keFZCuLsfmKeNc2V4/TvX3xZ8X
cpHeJ1JYv0qYi72b2IHTMHwyz1ouTg9xY/xLenSvE7J3irs5dGYPd9A02T65ilI+ePcIALx/5oF5
6vMRQo/XDjQqbbNvTS0InKQklz7IhSERlfZE/eSD9oi0HV7wsv8+3F2MvU/iAGod0iGuFfe5Wvbt
LGurQmcVJrIr8S5t18o4jZIucHzrCpi3vsDUZWf6qMf3iloIXFK6t2eFSaDSCL5jo2X2MM0P3h5j
q6w8sZ6hdt0P9c3voKlppR/qXsJAUJ8eFi1iAn+h64pOhWP0tBqG3DE9uLeCQ1+j+CinQ2zmFD6/
SAQVHcr3/N0o7JmhrA6lmI3oAuG0SueS91Uw4WWYh2q6H5Dmk7PqEGidGb5otOSy7VWv7cRn+ZT5
e0gFJz6ihsN4wUULYdRZClHp/lkKNc1bj83vBMgKhUmRgZL0ZC63J7ybwkB4TAJ2DTIrIfIrMZJ8
DKl/KdFJiwjSRPX4atqg+Ar9ONcbTVHGtIU7XDVZCKV6AyIyojWkge2YuANWgeIYjUOK+lyCCtbc
biNsvduX3ohQqkmlm8oWzLolF6sUlEws3jqfSsXkLszS4yemwzeg2tjCWvA0q6tqgPNIz6PnuX1/
7zhq8gAmKR4TWzhBvdzZQyeOIEjZ59MZYmU7AjYlzAbPUAoKTGLmKSYRx1pqrSFHTSBzQkfRc46/
E9OXbIY9yMJh6AqI5zTCbdga0K0tcrdoWqemI5M3YUzcSuX8G32wuSBvLRpZy3nayDBJLNkt6Ki3
A3m4HVYkixbzX2B2jZVbU7cSPVPcc6RtcLGXYpRi+ccbb5OX1lNSH8jyPhk3RxloQ59WkdVYvGlV
cpj0E0R9QKA57R4cuTClx9p2CkpsSaX3pFC7lThJ/5t56zwFt5yJMkHdoXaZeESPhlkrIS4nNG5J
7pjV4ocMy0kN0TxJB4lRZBWiLiX9P9AIsxOqqE5zvvRRrOicNzYPYLDRWaaIBf1KuHBKzgPXdW3a
Li5tQukUDCaanheQsG+AZMnHoV+Pscn+y9HifFQBCNTkkmG85yNERfLYDBjxVBTR8GPjbRMLjXYN
M1KqUQ8S0m0FO3oMySp3X1K+01tV44DSzdR3P9sy7+BUSUkrzq0ramEtabtTcDCm7lWByh99FbxE
+Ei0LbHUFtHoCoya4+zfUwoWkTBEzGww5S7HFApW9+AnY1eZ/r5TG4EdpdGsUL3BFZnjVsgy/Wna
oYL7MXZDaya+rJy9bb+CyJRLghm8rdffD0G0D1TM9MUsQxxq44gIzC2vRvSbggAypiZ43ArkHKXF
ZsmYuda8OD3+4guhErtIrAIf3KkDLA4pt0lM8q0QaZd6CyYTKmKUPbGD2TBoM1pSsKSJWPnYA6M1
BZ2CPPfkOKN7FTgoa5jh0W8kP3rWMbFnaP4gi6GDHRr0s0ZE4AG0AU+TngHSyVoztZyi5Agq1uJh
ls6tHlL+IBGV9SEmyGEvDz1LF60lyIyQ8K/NtdRO7Fkltm4qza6V6a6fgY2Bfva9XVm3g1Xi4yaF
xcRbDeKHqvo7pVbY2D2R+3o2w7oDzTUWeRozDeqGiwBDJo8zATCZxggMNIGXftD2OW8f8r4jCyfO
88XX4xzmGKcY0Is/d4paAtl+qdMgbC3fM6knJ4BW9XdrLanYWyPQbCnUmNlTzy0NrVl+BPNbUkrM
2f4TY/hHLdlcOwReUY0TuGi0SNo8/AeXM0Jogd6YNhm9N20iGAu9323V968d1KSz31IPIuSdbt7Z
zRgVE2RMfoLhXA0urVtBucNnBPSg846/fpUgUT44lEbSOdeKlNFJASWN3Clxgmm89j4owfzF7q7d
w9B0TS+gRHOmLAwDhXXAF0abiS6najG6aYQnITgkSQ1YA9uwOALgn2C7wg4LmbmTSbI7GI4/0OHu
qwvgnUdEGhXVk9M3ELA71x5TiJrOUiTOvBZY/btiBRP058aPPdDa63h5igMosLPfn4d9nX9GnrJB
1jAlqY2GzwNfR7labXwthvefcPcHxItcX2s91G1T1Z1Xe0rvxa85DV4KB/nxHCAzIqAWI66geXnR
8B/Kz3c6cnv1clzy1xR9ipNebGsbvFieU7vXTzRSiF+7qevdssEXcdMJM4lDSgOxsynHWzeTMa1x
FiWudNyUSv6Im/mpd4Q2KiwL4OyKmHlrp2XSmIGIQUR47SopcgsP02rhvF3aJJXo9VPA19cOXqp0
3CfkhKAKRIfzvAfcdQMxuGgbjr63k32BEWhEym0A38RIsrDNw3Bnqax//ChFGsIJREYMxvXAqilt
5DQ40v71oCDOOzR5H6rNlopU44i9HiCJFz/W47nyauUMJgYcIOEZivM1MPDbJ/zYAQ/3E2vuhrSR
LbJgYn5OJnYvefA0Xj863CVyTOweUJDH61O18u00GAHNh9st62qZbMoouX/sA5H6cCspc6JH7ZXW
Z6nTL27wXpduN16nso87NJIMWFcG3XjFzde1PyHW9ThYQgLgAIgIbSHQfPWCOmzVuDhleCCaIyXv
1YHKr9MpJ7eFz1MTokZuIG+6tTVI3Skp6HrKsxs/TgrajOMdSbI4RJIES5KkcPShkly6xNLL1fdl
O7bN6GBgd6rzSz0e8n6Ql446Rqc/ha4dh2X+taWVRssLI4oFY5ispMLwW7o+0sx2XvujwpDOn7yB
nDZ5dMxYAP7v8By2eZOCvwYSPgrMj+dDxV1XqHdlRu/rk4SX8oGHvxtWzuOwfIMvZshvaV+sXmTB
SzPvbbhxNy7WV766Fmfp/qwqLD41qQFUjIIgnIQugxL2G07YP3opuHqEB4CT1esOpuPbJJbE43N8
q2/ypnuScsULqdYbaF4yykaC+Flfie0XjuMYsm+eiXOP7roTS2P5WRC+12T0pcrFfP2iW1KkpHjD
kjdBgX7MpsF3P7y2XMU4UFmqC+zlKj0PvZZ/9hTWxzX8uBAoSGdO+bBp926gts9ps5sqnvU1TgCM
Hxo/1OSp+JXkPZQJIb0ZdN1ZygX8exo6uNgj+ifmbewkBHGQGTVzwmyNHFJr9DLI9vcIw3UwkWz8
aq5LPnhlKAhM/b/GeHbQ+REISP48FZi8rolC/IYkPgXXe31Hs0rNAcDijRd2/yvyscJANiXSVyld
An3YVskrhvrecSYrjfvZaTJoHUYN738wzc1J5ZjZTD+pgzlit1d4eTBGxuIzJpBrwRsn199h4f7h
LfhhwkHtKTn7JMuwt2f5qnOhXjZwYY/sVRiA4/4yoPB6RHUCt6HifZsvtCs/L0qUXSHys25C6mRY
IjSX5zqDyhRGjLACVSdkeyac1Nw/H/S6vTrKeh3vNlQ4kdMuNym04cfPrKvVjirm8ZZfSMKZmmWJ
8gQ0yf5RFuYSZtfmv0B9BbB+3ISuxAfk88wifqcuo10853JA68DDjNzvoNoqV8FuUDlfS/hWVaHB
9m4+2CViMFvmi7yji+MpTTlArzaDfZaC6DogaGgy0zGHzN5Q5DrUM4pbU/pnBeoHQb7DLMFuyb+a
EXLD14Eu+2V6bbAR0TfsA6aDa6A0sn7b4tkkVU98hvqi3LsdbKwhzHfWFRJiqnEg/dPd5xXK9oP5
lzvD46zBbSZJ7PzGyuH0M6zA56fzynidmI8ynQXG8qR7X15P5wovQ316QfCX+6AXOfVYcx2AHOIj
J0j/37+z6sEjwa9PUhb1zSc8xFORgk6giViAwO6QbVVMwaN/o545ukDfLStqs8KiKMfTBYQZguLX
bvq3C/TbvLUMn9WO9zCHlkhB/u0fKjvFeW8SG7HN5pLjq+2ezJbMAWz56Vb/dno/7vhWXHPSG1Re
tenUKHFdtqAER29SeNfDSl/iFoOSAcFAoviAyNUyBCZc3uHlB+NXHulY3qVDFqaAjb8othAf9c1W
7RouFKo6Bo2Mbet3NPVooBVC3RnBs4nqoGVHMJUZBg0InkiJElBF8qr4nTwCZV7sYzwTfkZ3641X
R2Wc/fWXziPPetkqeSMwH8J3nU+XWmPsOWr9F8o4rSaJ3uetAy3/YMpZbdD0cp749vaaqINbxR/h
CP8+q+/p5XeVJzaAyLDWRKWxZBHE9e3+5Yg9CKhPNalYFoOR8n5DI3ylPIJ5OxT5KhitJYuk/+hD
Ub24MGZCYmpLFi3Q6807qI2T/jb0uEI5iVInBzz8bUSaMDfCg2sqA0KczV6GDdStkbSpeoo61AGo
FWfnPpL5ksw4Zcg1KjRQsncuPLACJJq18z39VWAFZPG/SJiS5yo6uOf63Acdhc/6fcd6FoDpyuK+
GKxD7BILWNaUNmt0grzZvfjTUh3gbGZtKluLM2re834jkCWnoU0uRH3wnmoAN8R5y7VakDSJKHvW
0nSmYCi2MArovCMvjH/cwMofP2hF8CYeoifDMTE5o/L/oI4vg1aQaAvrUeq0KOZDJiiVk1YC/nVC
tmC9lmrVCUiwIpsua26V6tuKbwsA8T1h+iw+XUi1weKcBqHzJLadt2yODeUk2G5I5VSqN0iGXvKp
2tlKdEx6QnypLrQJga9JcWwXGWj5QXPwCYu/gArzo0LT0tOnzl876b6aQDEueUpJ1jM98xi/F78z
rvwSHRwyJlAxFn5cfsdaI3jOXQWy++XDOV+rGeDGW0NWOEEnLUKF3lhvyqntmQPperJXvgahL93S
Cq/4DaTp0i07Mn+SNdy96DM9O+QZ9Zc+qscsORY5H07BrZACOR9GrxvKsIHGBbnIsNMfTwnYkd9z
AycMQqZFNaW61L3MwzhQE19LyZqOFJnI5B0P6TrSFgsSlPD0+A08KINTTj6yUnQLi2g1evBz/jq/
3Kpm4QyJuk4QahDj1x483I5igoSZejJNx0f3dfEaXAnOo6PYvq9ehNHjxjAo/qhEMt5rEFRJzHgg
KqYSsIZIavMaXRRAds47/YSMmqyvN9liXd5AnL0kWxWXBq3XgwqMViZ31QtjZFhZmc2S+jPw3ou0
EOM//48SBj1UCnycWMMR2yf1NRG0DRdFzflk4gilKXq4oDpV/mbgL+4ovt1TT0rnQJKWzQNOczwz
dJlEXWPKgssa97pahw8UgIbu+LVIgVFpH6YKuCsKIl+3mG0Rru5aUnAQyLFPp3hkig8/evLSzC53
j4BIZQD7nF8hZk5mpH2mrP+nC7JVlSp3nHzy3TDVqTYszDdgZOu64E59kiYxfmhdFrCHiD9wSdwd
R/KC1nNNOuGawsZl2DT6U+lWUqLptgLxMfPrnjxuMny07auOuSHi5TZdV7kdOHtP6lJ0883vfME3
I+qFqcA0eCDTlIyMlhpuTKRXPxCfvOx7qO/WeT36MI7Zy8s/3hl62uFc3InBHebzg6yMYr5qVIOH
MykbXZT1o4CQx0MaP175ZhNVMzEQuL7xuyQFUuKabquMelCbxoVjmY9sBlKqTilMFnwyc7VHTZ1t
FX1H5BSSW7LAgtSjgXfT4sysK0d1sXbPBLIdo/b4QE7Dr0N+PTBI69C/Eds+iX/1P2rerG8uKuOA
ZfEV+wwQTH27e6McTsmUma/5b44Yc7a1wN5dvc3yCRtDLr6w2qMYIXvtLoLekfTGmYmyzlrRR7bR
g0GRrSgvZFhM0ky0YXHJ9WQNwh5eSgAY33vek+pz7w4CQw4zt8oYC8MzN55pz4AC2BLk6/uXWP7n
h8ZPbPBxVHQGQKQMkK//SyOv5H++0wddjE4aWv+GF1Lj/GadHeXoBKSznm5cMuTVxUwMHBIkyBsb
Oqb6ykevKd6d3Hegxg+dKPOaWAJm3IQ2jgUqEyej0W4DqpquFIEPDfqYoM6Bm4MLAADYXnxKd1zV
JPXA95CmPr6MMWkRPOaAr8wSQj/ArVX583e2xFAocllQE6qvISoCbFDtSgtJ1GjC1hegZcHwQcJ2
fNQGmrve4JmKmNclZYUTrtTRlHBQTBEdfx/jznskFATyjsfQw4hYQcGZGiQ3l2NNK6Yt7h9+vhI1
U1bG4lU1trky+llWD5juvdkfG3o8OG/sSf4ecqVFbzlSdHpGwaIkh9GrPF2Ot4Jr/yFaDbr2oygu
KTl8hsxzAvCbcz0CloboZ6Qqevx20x22vS5QTuSZOO7RmXclzNYVMQRr999DZgjVNgT0E3djbqFO
GXlH49jaF0f+T8W5qDKKHAXr/5PDcfGEMZIi07zIKJuZ91UIvn89vx3B/26KZB0UNEEXmy4ASOb8
5LBKthPSE+lgyiYyMzbmFgi7pUcEXca0WFBQvr8dAkvoMi2wLHALduQFu2NElof2s+gyGD62muOi
0B6BqfKP0iK8yvfGSUJEuLmG+V9doU9zPZLL3QVAPCUNGTGIrL+yjf2D0Bt20rpPWNGYTLvQQOZn
3BpFF+4WPRyA/0rTDyrYJiK2+Ysz2BKd3EGT2Whi2EfTxs5wx2w6e2NB/IttiqYZPLDH06QrhQYL
EqQywzdphJn7xFSG99kB6SvrYzLRPGtdjXwA9mZUnSPHkx4YtsodiFGSbBfEy8CSow5nzFERV7Kh
m8cWvuhRcV9xddzRGXJjdLahiEOKLZciZ2rouLek3ghXTvdb+SyWCWsmkNx5fEoHsc++wMczf/fO
wjfNScof9Yka418ITOUnSb31Gt6VGTrVWTwMchzS7fDXrYF/SupT3tjvQmA2ShdrB0lU1KBT6IeI
EJouslEeblf1ZugKIpuektANC3CmH8YtSW0Vj/b3tSCY07JzRlW6P6BP35IY3g3rIbILWnqld0L3
qdgH8Yngg16HT6xjthnOgUXPMwAAXRJgKDAM+BcDw2kE0Z3NvVYihsuxrByFAs22UmgNtXVEnWm8
1mKoplb4VsQNQd7oQM2PYgzTn421Z136zGwjT3T3ouy4g9Xz2WEKoM9X3VHVmMGibabIV/MOpJTN
biDbdhH8WiqcJ9PZfgGwYmzd8ziWiNI5rbFayK5rt+prdrbTcScaWwuAiPJdDNDtWxDasA84wtwE
8dRfLE0OTsN60IUUx9WUx0UieBX5E+bd8Yk7O51VEBx6u4IoC7aqbwd56zr0Y3Gldf9vdNe+RaOb
DJ9SDxm7c8Jm9gg7OKL2rE1GwdedxhFIk1CuC6i1QT/C4zZkquAPJ4UX1iuuzJoDX5jaIUgwPVbY
EPEo0RLlFEUHo7MyD+H6Jxwt8kFGZg8mHZduwYCwrJzn8HNIVo1c3fem3NAunsrb+cpavhlIzeIi
do9zSkX1nbK50W8y36OKnzLZLi8aL/WnN8w3xMBNggacT7dHLXMMfFiDvjLgNIwfisMfHVU7jA7U
rQGv8+PWB68cbT7hne8FGz7acXsW5/ZP+74T6YsMwqriwssilWtn+0mMTLJLEjME6mfebeXX419n
QiTWtJ+xw8ueJSf9hM3HPWfBxvmSidK9EUEh9/h3GaasHV58rIKwAdDvB5PtWlwUivI6v4jYwnhK
TxaujZ4TJoJvqZL3EsYTdj7tdFWddj2oEzrqHg6JCjIfn8E1axWF/Zmf6CmEkJIAg4M+4nhleraq
Zsj0EjjKkEZgPjq5Z37x8pnhRgXs/W/KpyEaLmmjU4Hvk9j3A57CvKSr+WpWrz2AEqa9PnPWkLji
MT5FGaasE4ZPGzUfopJdk1o84wLWtWTpepEIgCJh/Hd+5lOQbIqJZuih6QPD9fKfuLOmUiwH8Fc6
x28HkOYiqNqtvO+wtvZPxdWjTzZbQOPylG+SqTNXhK3LhI/0Kgy1DlzCa3UREKDcPKVUQ7jzdDlK
aox/NO43muTfvQ5X7qdc2Ra5/kk8BMt67iXWtjI/+u9HdBrppESjNDUeBRZyfaT5ZnT5dyPrVVkM
gX4f72Q4ZmYkb4/wSNdKJ6L4fA6jG7QrSxfdMkEgWuSUgwrlm2esn8+yN589hoKf7ETb4MsRtL7w
qEKGONAwFGiWalTXjnN+QoNQ8QeREeC1Hd8XfYKkBGLCkbsFbeZXtwoS90vQIUogF0xAeBtVPBei
8Fh6MP9SheMbgXuyHYK/OKSayDLYM2/KjdWQQ3PCIj7NRda519VhZc7WcMZx710JkVGHFeEFsIHM
u0kZLFqUD/eDOH7hk7JOO1OcyyBYmmd0EyqLmLgUC1/BXb5UBwY/oX0EThmGcm+vWRA3yfMANmQG
Bb7dtzees6o7a2cOPPMHLjQ1RqODvAPGWtiLL8/yC9YeWW61s2nscmZsI11tWmvhgfJvOv2X4l1A
DS35XvEKpAN+y1P0lvY6ABP7/XOcPb7REYRFI+VkiXyBnvbMl9AbycSdXrzmjjYz/ZsXVrhRcn8W
WA6dc81y+ACkL5o/xHHjw69IHCWQmAOM2d2lakOqEcF9Sak94LT/L02/bp8ELkjzfJD5XbrdzroL
q++LO0akiljidKRryEuZZI/KD844CaogS3GZ8JoGq9s/t5i8baX2oDE32PqNew5sbcJT9YTpaGpN
w44EEjEpjCrVDZ8RTgXwzJ+iGnk0QsSC9jm1YFnzMEn2eo/wzax288m3tZomhU47bmii/QSm5J7o
vylS4bN0Kkv79lKABeXbJFz5JWsPfkf+mQEXhxdJeGs2CoZbdkSab8gICekhkEDu/G8A8tI/vEt+
yeRZVeRymAVyXappvDT91KnroIMGXgA3Uzx0xmiAxiSaFx+osMG1tUup7cvhc0ucpSAIp8D7jk1B
k1Ek3kMVs6lV/EB4+PNXrpvIGx0PAtgIRpsG4HWFOwy9lba6EEiibJleRifOrLa5GndhCvi4CQ30
3kDTmXn3F61hftUC3iHBM8v3XNm/u7PnqQef2aI6JdgvVOWOaHcB4jvHvobeyETyYtYjn6MJFHng
ePwIuH65XI4Cr4hGPy95OU+miNPkc9wbaJP6brlHl9eI9TGXQHG6rE0bJfa6581fVH9Si6KhanGO
Hd7VX2Gz3DMD1OeKvGrtC3xMvRylAWaIZU0ufMNX2fvj4wXmRMOVo4SmQzSme1QOLgd/oKHggA7h
Y7gQdxlgge39dtD8ojvMnv0iEFxM+svsmLwMwpyVOjTfTyDjIVDeFTYRuOcmR0MiDcxlMlvJyJhe
M0VQlHbUj00H+FYIBitQjsg1ks4KluOxlq0ZAxkvKaD0LX5bUUq4bKlgcICzAA/K16BGhwGflYdl
AJNZ8h1cWMhGS4pe3Ptw5ABhf8Dat0+Q/lkOeRZ6mD8gvnyqLUh9XdjZAxEMmnVOhflwAMYvDTGJ
cB4pdglrTbU4Rl10ilxX9DhiybxwlS4ayPQ4kOAF4B1i7wMaFaI5Z94dnwamZCRyMxNj4eGuY76J
4D2oNMMc8FSyytOKpkWatWtQyZQ1CA/jm2w7/pOhj7zI4L7bss8FKrC/VhmpJAJAKOU0PcW+JXtU
Nz7T/10gvoaoo6SQJQGJM3XNNPrN7jtKkF2dgE6Cyy63oxQdsWHZTfjVa76+JO9Fw7gfqG8Vk1VD
+AJADe21N4dJ6WD0izBfcjqaHJSPKo8n9mLxfyDyeU9vYek9dWYyFuYvnNAoFtmaENSzBQRs1utx
ijNDLrkJEVEk0vYYJwB9PrrizXk3Ewai8kCSBahgmLSYhBmJL5Q82Pu7EMSwzKhZ6wlVdM1JAFQk
/XgQ/EFjdUQRH/2Ni5AgVG1Fr3RGm7zl1zIe0AvvifnKiFEjL+SXf2brqHw+MnFhN8R6e6qpLyJO
2Wom7wo1vHkSGmYcEfEB8grbg3B90iPNqsgpoNzNNEWpZb9u3yEbUOcrHKGFG7WX07S9DLnYBhxW
4MuGCBbu4Gror9+c3yNl7oDar7sfTTYBKFVkZSxE4QU77O5f5AxX9z7fNMUgRzGnIbw7oMBI9UFT
iocL4wKF2VC/NJ4kz3ygoNAfyVrtwF/Eq17KCKFhpKorVF4z0iqz1Ip08an5NR9EZGFUw3JLRlpR
F4emhBFFkAphMZvS5F4qAkCB4uQ+hoCSitJiHsweIt1RNQkBVdjO3P1E4tGiaDc2Jpv6U89iUPBd
HBEITcOPBfb2p42o8/Y6Q1B+rDpOpypwRIljxtDrnYufcnreT1DQdrtcIrsnh2aa7Qud4FWFIPkX
aQyGCQrkxaUN+kohowmOA8C97zZspuos/6u3Qfwgw4QdL07X5hfrVVk+/SVAq2bGLy1BB74W1SDz
T/MhZhcA0LttqfQZ4rUEnXOrra5nUbd3+Rkq8Z3mZ7a6Ps8yfGR28Mrm5iVBU573Uf0Yf36CiHqX
ATyoE8+E6wUiWCYjSJ/LpGX+KL3ihKSNOVX8jiOkDrS00r1EnPzb9cAdWuYcZpfygzxztO+9QKDf
ZrvFqsSbAbHeMHfXAURCReOg7d5ykICFp+GKvK9oJD6ItzLrTV6WyFgsJIVywR/WHW0NKhzZw4bQ
amB8gQwdbunBG7Sh2aEA0IfUqpHi04vX8anE5hes3cxrhkOfHGpo9NP+DCF+51UdX9KGCIDNFJD5
fxQ7WxUcYvN/xT5QcxRa4RQIScc6zgVbL2vJ/ADHKJNPBzPXrWDaGC6gw+yQpW85AfLKFeMjRlDh
wco6caePbEXQw4qHkqPs+I+ogkYcx4MXS5tcJZvmHowwLYZSS/RhqM0TTad39rRr57JtX0hfH6iD
wJI3U7lNJH20OmiAw/YUTkXHZYR4dvuYfap8vnqk9rs3sun+mIl4F1DHLu58PBskVWOBThnpmz/y
na2fZrI3gwA5KFMDWEngBgNy/WH052J7TOvN1bcQsWRxrQf3afCP1cMH9dUK7L0Mluj9wLY2yRp+
kR2ie1WKKY2AN4Z9F+9NXDI+U4RFRjfqX2QfX49Nrv4323PbI0I1wH9T8XG0VUdUHL3wxPST++X4
dw5o52Cx9zJTLasnPO7fMsBU5YBK/wlYO1exSREmerVirdovene4xlnQZQldMqXV3lCCGPSkukdT
IID/b9DUmy5jTV+4qkxU7BgjZM3y2e8N4V3edGhqd2MvL6cb3TG4oVHKaAXu4Vk+HHBoPFzCmjY7
4I1+5fTYzOSNlMa2mf9zDe6L03Ziw5Vud15XG9jC8Waw7iyFKhPsqhAGlk6zCThuaMhIbOJsQWff
MXlZZ+o8ksB4GATJj2DaI61WgOMhGA8fqQdy2VytBGWRrGLvKbVZtIw6Dvm3ilXSc4KCeQOEuiVl
6xSv7jN5wkPav3FFdJWV5/i2a+PPJtScSu8YbIAjVVu2wGXsls1fqfyUZMsIEpV3OIsqiOWt9O4v
uay9oZpV0est03OHnogPdwXhiPJu8ATWhccTt5EDOTg41X/6I+FH4SST7yCHgj/4PGEom5Gj07cV
Uz5x+z9jouV1jWcIYFfjvajgQ3fQzeGFuNEn+FZkIhNxybsVhOnR9SUHpvmCG2u9LIZxy+LolTLC
veKLl+M6zuJqJLHl3bVz0X4IXpCJ8z7wYVNzBeBm3kKRCyYACYGV8HeGcPFHtI5eaw5eTdybvcPI
7tmHYdMCCj1oFLMwQailtOzgjkvmRQb+GZgi7kWf5ooTBECgRbjNm+aa/O63xZLU+vxJ7vmaUiW5
dtrXUe0RWXhDTRyZtMG35kaVj+50Gv7f2J4VLi0ZLMdW3oDBAFAKUQyPbT9sjC5SI0NbaAxfvbBQ
gO+5zYHtkOPEW4mUoPGzjryNduSmhMjGbxFhAS7Tw+rXhutEoXj8jDukFzABzAjBmllCf+OXNSx9
M7Dkr7R9T5odRDwbnAdmcg74Huj3WsTSQpJx7lXhe64o9/0SArgMF8CyFkWKRoNpCZekGAYUpKmN
SX+xaDKa5DI8rlp7SoZhZ0YQv+mK2x+9BVmWabXlInSewpLYKMpJwDjIPYD144mdHaUe3UJjW7xX
OmB5UVCkxr0uO8djNrprYTf39mGm/wAFklpxMHO3BqkdkwNlQtbcRe5cq4v7pH/PPVD7u/XgwjEv
1tZIGsRnUjlcSJVWmp1iEiYl6Q7odXVgrFevO18MYkRK0aY8pmTQcA53CPDEcCo3WeFTgJR2nVp8
ZCdu+b8e9u0GDNzyz6JmRyYqhbP0a3bmxSsSwT8GTWrlkJKbb5flreWrVze3Hhaxpu7wndEyVCG4
+mQukM3vI1skmLX7o2M1HckSMTJR+Ew+xckMEhFROs9Rc4Y78t8AFhSvqnx5qismB1ivzO8izHye
KU2vR1Jrd1zdUTN1xjIZo+GNF3+2d+pKniWC9aN5/5Tf5oli3MrLASzXFctmF79vBeL8SjDot0bb
mZr0JyIQsXZJa9T5qPKzoBpZDMzPozNPxchS4VBi20Q+GkdKQL0jJunRR5z45IOT/hug/JJ3NBOD
NcDLPkBRajAOPHkVZooGW/udC0ifVNflapZRcJTzL1H/bBZJ+uxZ/zOK82+0Z1nnU7+LmvmygO4u
xwHim+RJe3JGeL3vt7YW/ZS5rQDiV52sGDqx4x3vyAjcdoB5PDG40+sI61AsB745kpLzYEe1RID0
A4Qi3bYCBGGxF4yvIttR2WwAw9rWtJSVCE9cF95LtKADkE1BBUCTBZbA7OTCMzSOgvWePtC4KzSl
GAjqPz0AFscklTXfLMOUZ9haF8JA6KQ5592SxihZcFC+1ULMlfhtuP2XiYy/z6vAYoTY/1CPskrC
jz3k9eS9gKD+HFlazaRtWWOh9rNEbo3MZRDhypGQ3fWsdDSTwI//CAl3jf8XgX/hP05f53kFVLr0
d3PcakvOsAleS5tLNZTw019OVFUW1DTylnuC3EvYeMuYjJcRajQ3DyUqJ95bcRMt30CMRB9gjiDs
ZkmEWG0/JU62HXgReg0Uu6L8duDmXrv1jdgOEq/Jd9WTu8k1KOdWubllLd6UydC1KYTQ61armPgv
YrUfvEW2CoUY1X772SWlDji1kyrnwgCHCAjxMabuCw9Manw7el/HBpqGRqs/NdcAMfRwWD/GRPQh
AY1egLfzJ7ok3KQbtAvjKWkk+lQ9QZgWnYjX88r7KSCKVv7dvYqqdbikPzK4e4JXAWBUpfObkh6z
05JmhlKWvPBTVgKI3NvKpnblEr/HEM5junPIz+kAptmWro2YtufOL0NMhfP9iEpQ7W5w7LBlLzKQ
plrS5wMHEJVQ0U1vAZEl+VPjtNvbZ7G2ouHrz3Ddg5EqXehtgCIshJaW74PKH2OFJ5XNaBifqb0j
sNj5bsrrzWmv+lZmHOLa9KYsWCKPgdFLomRL8gQvYLXtPuZrz0Aey7ya+5JX+reKqLslLuHdq/kn
qtZwR4dLqkIkodoY5W45DRPMhgzYuWbrwZu9F1a7sso/mVw8t9jP5cUxtxWhrbtrNiEAo1Q44fWZ
P4qUjSdNMumDKo+xwrQMyaEQFJ/l1/kKwZ52DpmtS4eALqyfi+syJYw3oAHgqHT/aJR2qpnKr+/M
Z75ms3/UPEPm2NlAt4pYqC6Gfk5OEuP52uWGMf1Dmg1cCrwyqwPAwNKjNTmulGFRb4W4OVUyFVz8
ClhpLghbnCWv81xcROs6CHO9n3sjVAlK+fqwk/mIO39l8WxKDEgTkQ88IBrDzqy0QebEHOZRe/M+
AvZTe5cSVjfnARqkvSOPkndbBanOhx4cUVw8FkY0IZiZQ0OgCzQIpou28sRNWpWO2YYKmJFMiUwP
D7MhZI9p76SXvwyo7HlFXKG61RKDuhBxwlwlzkZn8IXJN4gRLv0vXxQPqVoW0ehUWPlfzi47ev5x
Epc/4Z8qMNHShDTcNlIWXN6s6XWFrF5U0NFLfpM8vZU9LPkEnVoxuBU3TKQ3lZNPZQ6OwinRYUTd
CfLnajHbtUxZg7wmHkWp4TkFl3vdRxdmdxEFOwku6PiG24ueixI0Io2jj1yS8WrHImMxLnL1IpFj
PObAo1c5frGwvEnXVHGdkRgIIedg5LWmIwbwVhEs+O0nxAeaqRiXqw8kHb9qbso8NVbeJ1riSQ46
2Xgp4Vc7UjME/x5JkxTcelATZs7SJDtXJ2QbZOBJq+3lK53cJ0Ud7r2JhJt+/3ncAFQiouqCjz0J
JnDLl0uHVmlZdNcQmptFk/sEFN7J5OQlCHJ1SysKLp2QbXBUieONBgTv7/t6aEsWmQfQRNnBRMik
G7Ocj3UYe3MsyL1f+79bFb52SuKvLS1h8ndZFINJKYlT1AzsCUYpmJxK6TQv0w1A1gakX1BQc+EO
qevPvgA9pi2M3TrZUs/gMcEkiqq7OpLonU1hDhL3IV9eju7VNAJgbG5DiOlAcv/ine3C5I5Wqu2N
vSb96t88J4MCcTbIQnSJVBlldUcBaOSsh7QKYEEUQGR4WQtC/F2C0FyPLc/9R6c+T8u3KHoZwcko
D4xzVsiYyUuNJSjgNOtPXOD90+zZI54SDxk1uwvu5Zjgc7NKBrmUx8HPlbabtLo2PmJ9NBKf7LKU
3ECRVkoh4ASCl5K5VFzRaGMUTFl4Y8n0pGp4R93fPMHRDWCBkvUZLCyFgOYZsrZORZ1E3a/oh9tq
q0d3Yvxf6r6nhhqDiTj+W4HycQmLwD53mkkBjTnT1WXB0Xn2mlDsfqxoqU6zViQrRDBnO0CKw86w
ELFpJ92VVPLMa6r+CP6518irNrrLphLZhkXPHP+4mR+ype1nEhUIHs5Ckg5ta/e2bSC343jMMfEA
pVt3NO6fnQ30XKFUL99vKnxB4U0VOp0pLw4PzUU4WENQ1LPixRV6MYGM5Uw5C3nTFnnLCfI5SKRk
W9J8B9B1p5F0scsA7vMZW8SA/Z+bTRKGIA/BZ4ESTT1vPTq3ZRJ3wCCVu+StO/OkTHxEka4KxwhQ
mwsFDhJNmODiRPocR+1foFDNmgs501BCtBuIQ/E/wi3+nxUi23aoonQUtteHOcNdVxNcsMERCh7r
xxQLS6jCBvAggjpL4SSSq3+z/el9X9S82s0Gua89Uj3J0wMU+Qs6MVe2YetHXmQqfVFmSnYTwUKa
Bf96YOpUJkP8lqg+0AMd4waAY8YhUln6zZLpAYQd0Fzg/juoL80Rz9jNHpwGyq6pJ7w9LhqX3vGP
BQjmwaI50NbEtQLVs1YJhY5OsFov4QABd7lD/Crf+zZYzQJjwJzJqr1wDR9yJCAkp7zmqElgbb3x
CXDmJqD8OVR1XZc7NMXW53U2lNM56roR3QRGRvANZa5Zrf5bhWFRGCX7PIfAcJtj3Z9crD5qCTa4
bBGusSI4GSnop9kKJoYQlETLH21KWypLqUFHd4rWzjniC1giUbz/V3ehKNPwKZEu0MKy6Qt5Ydn1
FhKY2oY3GJx4F9w292vGDEMflre8q057DUavgMqBMas6Pfx3monAzFWM/1orXR/4ytWI3bJhEZOb
Q+noajsTeMvn/2Qd1tpL2aSNu7bE8ze1Qx2X+UoTPf7zzn5bGlCCyiywuddRO0mKLX2qaYOT6VN/
KeCDbhJ8P/jXw3xaWCbZv01qeNJUPoDmVUXgdUHYz1y6PJSKzndQYsOVKTvmjy9DMr3YfNgI3f3G
YX6LaTIMMw4SHyXy40mhDP9yEUCI3ddPKvW9blqNieob+rWWl5BZqGJZnWzns6t3PxWzQoWwV75p
ofaDPvQTbU0c0FgeJw6nJqt+pR1RoYrW2JAwdQiVCKy6DUTiakITlrhNJrDUdSEp1EzurGLqFTqX
uSLRZRUBLFC53urqdBlC4GClo6LLqRj3cJURGpra4NlNHITgJn61l5q+kyMSBOy4TE4HP1ezJyJL
thlKbMviufnjnisVDNrb5tE8G/AE4ZZVphQJt9fkhDRrTVwKWeqtlP23eTHKuPTFdkPUwn8RNM+Z
V35eCnL/h5lN0znPjO8tmUtKZNoWcI3+qVutzgQpqyyBarfOkytQgAY90Oa8cxScWV0KfR8X44l7
LQ6q6poXnUXeqL2Z4Hk1h/0o13snx0YUmKRg0cfV/DyRntd/UdR4kPkN5nCIg59Whkbc0l8Oze8j
3lQYdQM+f56oXIKg4TbOkhYDBQdI+0JGb2dmC2xnYtEKn4NErrkKOhJbtGkEGAgmghu2NuB6C+BV
mXuQNRmAJzEwqMHPnxPvmKI3zg804hHBTmvqaUETw6Iuz3DUzIRZBeDeVkIemrw6VAVIUrWD6FYm
06lZk8Abr7+hTur/jd1HRn3N4iS2/LH91ZIPDUB/XKAPD7C5EXbJTG1f0tfV4jQju0lc6Y7joKNp
hlslFisafqRK2zg7PHynytIkxJkF1cJenqL0OR4MSuvyEbIMBgweG2kgrixnHClJsLEI5nEP/mJm
vEPdnJqDiUiJnM/t85rL2WsNzMyKFacMa+VD/9azf5/sPl9yTn9NGWHUvJByDS0xmjiuCdMf/VIk
5KjyQLIGQSXxjWDrI2BCeT1dCBTEHjGSqgN2rPJYcLlUhQ1PQnsfM/7Z4LC49DCCDHFSTInuiuqg
aTj0Ku4jsHXVi9J6b7EKMf8NLSbKGY0o2cFR+Cy5RAcC2dGCCIqBJb+Uyu3N+dzBVbXv9qULxDt7
JDzszbBIUqHbFj35Cdjh2Q6qNIX0hRJZKL+mb6GVjK9JY+Y581alZ82VwfKyp88NavkBjDFTjiWx
BiegGbO8hYtcnQF5aYmGPzXB2FgJKO7AuQS67NBaICVtWVL+2nq5Upbbh0ufUjw1Q3Ob2iWbluFT
gFCuXvW1gEW5zOhCihLqhw8oZCQfH8a1hMwWIduDYrctV2WKIe2iEIGnYW9wD2/w+rpceLhEz7za
Ae3HcDiK289XzQcmXBryEcHdiNr6dSkm9043hdhcWPxVc8tm4L8CCUg/EFNY1vWJJtt8yWCwJLTn
GWz5CnC69P+G281dW48DJAk4/Or5aObe2F3VWcfTIPfSIAV5xp2v48RzUYUObaQx/YbnnAsZoYbp
hPpWGKIVuCzO3QCXGvqOYv+aCbH8MgnZElrrtUCjcedhWywFEjBvNURX9KJeUOt2X3JiVKzuCKlo
A/kLU7b7J/E3QiMZjQtvPeaF5zIy7iIUoJTPBb9hSe5gNW/vesSJBbYfRXySWk1aQISkYc6gkqKS
6W+f+BbrfRNRLB6IAU6jh4atwz7roTDzpXFhx/goYgauDE4nBxtDULZQiVppgnKoLePVvh8btcrB
xCcuR8Dvl5xxTSsYcqT07JN3kOZQvXsmHOIIbmtkSHgoUTirS6mERsqQYZXlTqyyxf9o6k65GN5o
Si+npc+61Sd5Czb0Eh88PR+qmhhAbH0I6WsakbZ3Is/EpPeqM9JN8j3c6Pmqs/0KDN18xv3EHkA7
0qBm+c/6eDQqLgH4FEsw/f6VQJEwptJ1ffdXQQXAFI0m0rWjmPtzAkPDf0+l2/nb79AG/ySndKXr
qj8fImajYzsuNahYUrFfiyC3ZftSya1CU41IPiaE55iuccQvW5gH0tDScwS8iBlSXMpEMNYtp/L6
kTeUkq0RzpSdxtLHSce5sITI2bmLpQEZxp++fDIeXKAiBHCuFkIe4ByQgJ6DBfhJdrs3+mySTYl2
0Qt0/T6JdanBhGNu+Ft7jGtdr0lUazLaiejp/+sSKdKrj8RHJVWalQvdI1l4a6zAQ9i1exsCBLUx
cHycDgz/e1LAH1uUSjhA0BBtU0D/IgDQwf1/fj+j2T0oEisl7/qfhWgEAAIOC7hV/Q03G5SFvI0V
/NukFdfmID3Hgks35/sqt8bklgYxG9gjN8VqmVXCj9D3lir3A1yOVGBidudCytrC1PfiGhvE1Ml0
+A266JNI+A30tb6DJt8OMPf1XTwYLM7cUiGNrsxSz9dKyXZ0YYw8KiHcM2oXv0wGpuWgMrMrqEFI
K9ZttA3k4YC7FgYZTzr/ankhdEVGgk1ygLT1NTlyelYsHcwjWzOdmRtcMN1d86oSXUQqgYcmlTJX
UbytmhcRZenuGUZSMdZLaIevNKXG7615WQjfyRC6ynRJRc5vX/eVC6R8wFS7gm2msDYMqtp1fIEd
YUSOCBT1yQ2T8Fd0pSgdBOTzuKkyqLy0Smb9ynaLeryMJ177D/XQIP67ablDP+Nx0axIjhQOJ4lr
U6XWDgrAb1g5iAydZUBXO4krZmNfjLkT9Gg3KkmeuDV5zDjsZX7m1LVtb7x8af5QSU8MjiMiroVx
OE4Kk70i8xJnTzjI+MxKRLhjJQvnlBgB00mdT0BqrwHaJ3Rxcj4kQbdRM+1rDVpZP0FnnGny2Sf6
uvvwvdXwHPPfB0oBR8F/vitcpmvFuAocJghQ4rre0QU0LspGTZcD9aZMUwcHgAbyv8hjEMWzOW9x
wnj3M5O7MOP+XfiqVjWHOhBHBvt81UD7rn/y5/L1WS39BjEeKUcLrv2ncCZuXset8qH1nDp1RaXg
eg1wHcS8hCKw1C5TU97mc8LGQ/jBj44rClt74JLHx1NuUOVaiGqWUiidDJ0ujiudd+K36sR9cIf9
3CUUl2cu9ehecLa2yyMp2RU6g4oqOxIGen3KkaYRDoOgvCeth7ZaKM0GDoeliUrP0AxyaGhdTXNm
VoF81W2aVgBXJ5wMAID39RqMlZFbEhFU+lk3xYjVcEXCZG8kOtLuOQ3KKdhBbltK3+L28XpFMVum
OMpJluAzExjcaP2cI+jUCdwdv+d1uzHXTE8meJN6vyy55n0h0S2rjpt1pVmdW+wyqKaSgsC59WEG
8dK4rDkoDGEagCfVm4mMGUjQgnUMDi797ZFd+u397zPo952WyDsTkG8c8j/zkESciDrAv0wGB2aK
wnZOPEYpSf0naAy79mug6kO97TcYw2o8qlhhtTYR3zEBbFkWgSI/yCZ5H13S40isZfsd8Bm6+co0
NTZwmBl9qXS/kulto2ex9ZtjX0mtTAcJ0YTufReBX0lpGlQwEFrYODgXban1oTnD3ntT7/kRtNXy
yI4oQv8uZqFkbi3AN6YI5/8uGSvXy4ebWTdO4JM87GnnmqTB60BUuhxV6Was9IfzKCW+tlAZnVti
9iGzRWP17EsXbm/VHOglTgUYNZ/69G/fO14QhzkmYK5ikUYYp64HMYTWdqPo3Cn+95fGN0XR9Qah
MrrTeBQgNI0nCcKD7o4RxwQzz6xZLmhhtThGRYlbQxas9QmEkHVNgy6uoCstYw5Tpq284jwLzink
JCTBzgtbF6XLxMJae2upkQyKAe48teIXbAO+pNjUDf9PcVnzsjYlhjLDcGdd2+yypl/DrDFVsz26
Ryg3ej7AAtzGXt3CWfkw80J5sr8SF/KcttN4s8UCJgdqxoASXLE2CtMI63SGjEYhgEIoBZVC2Jhp
9mgwf5VYbTjtayHuWxI2CF5gzd3WK72mg278LHpDyEPvqFUJCT88KvpWPFOEv98XW1Z9xrbl0JSk
QunvS7CSIxZPwn3Q8ErsNTRiTraFn0VOHPyTjJvl9adL3lX7NRQAR6vixDu7F3MPhZxuH++2aNRP
nNC1v5zPgQnfQnTTTj/pxWonMnFPLrcGbFp5BZo1cQCitUn97/4T1xenul/V6De6Qyp7kb+z5EiB
dK7xqT07u/xcnOSw9U+9BVgkUAXS8KFsWs1Q3ksFLl/pZsX4FIo7mVoEKjkyklsPsCw2CfZWeqAj
5WJwlg4MdHAIns5uirsfmh82SlNj0aHrjZMb6LFmlwlZ3L/R5UnzKeroiUMdrblJELNOX/KI1oLh
FtKuVZ2rMatFiMSaVjCjGUPtpadN84yAtOlO5aWmulK+m3c1uXMMbVNwDzZatvZxN2YZudxW10f7
9TTW7xEptLGvK4WOdxO7v2W6UkfMYBLRq4wFwqgPvV9bm36stenBXTCyjNivlq66zlwYLtqBiqXC
bTD2MQ1AiyAi9WR6fkj5SJZlBO4FJvQ36GOwGSJL/oq0em04GXQaJCGEXWMebL1TG0C5op5CUHCi
uZbFwWAMB9AW7LA/9mzICikQHBZXnfivAd/En+WOAs8ocOU6WcKVKSRTZTSpReZ+WEHeq98FJE6V
V4efygDZGxPAA7jrOC71pVdLmqkLD3i+s01lawFG0g21K+lSde+yAOm9qvsMPTqUnM0dQmbon+z/
ZNp3p0TtNFTqkRm+jbH0wPPrE7eMoPlys+zLW+Qd+Yd+2UsmwIwG68UiUbknES4gqGNSv9OMo2Vg
UrjTpiBfQJCf8MZFGGherJxP2iwiueW9zHTjyaCRxfDRhYPqLMViPD8YOhZFjfqDEjkws1fGlG6I
3AnH8YP8XEg7Ba5j/EATIUWv2AbQV21GMzJjpHF60dd9+vaOYMznvM4v52bEVijRt3z+NPtys29+
1U91kV7P8PcGg4SSdMxzfnbSfHrYTRmAGSOP5jsY06e/SwwLCyOQtuwGUe+sh6qVFrEXByhyXs7i
pKmswrNuRErYluBVx45E9hutXxjlUOxxCC7gVOateYimQ7VyTyMbKt1N1eZ9X0FZU8nLbFxmKwQU
4gSbe/i+Fvm/r0w4MewjGb8SGpigJ3zLqH3hQFTKKCdGwwO5NpQYj9QUnMM2m8z2KUY7MRzOLE88
M3GuunCaOcrZpNH8jxKKgrcgShLrP/rJ9eN93D7dVT0M3nQ2EnWGr3xtU8TxGRetjwyOKMqyMF5V
HZZm37Y3dikD7HxR6TUKeFZGsYMKo+ZLz480bXtNbY9rWmuVFlc6/NC5BmxSsMEHlAGcVbm26KAn
zmWYm9IxbDFM2ittv/pmk29NKpMQihlDooAQrHWqh0qOLEz1N8IBwRZJNo2aSi17pCtncasgae+0
hDs8OUAU58gm8ZCx7ixJJX1hRWB0OxXzsjYtReilsQzkhPltfjC/dVM5q28Or2nxNybd6mSFfFZs
ZuCmMsLoFVLM6M3KCF5pB5CQ5TvW4pBFWLXmksio3kUDfDoFkl0QtmakVihSowBngKwmT8CtZEPL
Xa8QDyMn/Ft1AtJqBWf5JA10taZzbdxTfSXI+JdyvMu/9OPMGkT1KvLNM8+y4Dul/kxFkvZFngtt
7jo7ypbSEgR3MHBRQlfjprIaI/8OkFvkGIIiTO8qBKlQoTnaOfhzyVyM4FzquXvIixN17vlpXwfe
qToYalvrAg2Ix0Nvju2COvQ2V8WPXvC/44w6sUAIv3EAULtKz1g8nl5IOMe/1152wdu1celqkDx7
OCVIrMT5mIUA3GoGD3XzvjHjm0X74m+v/RborV2yOaQE/4A5/LIkumeGEkPTlWa2QV7jryAlADAr
eMNDQBo4thBfFqsmEn+SQKXp/gGQ8BKE3Hc3uON/WlmuSiApTY6z4t3d6gjk5Gt9AjktZrQ2NBZC
gsmsSqq+CbtzTnmppuWetNuglTcjGQhCpm8lNIo7QPt34Ae+5gj8rj3m9gzOzKsHXzS13WgA/cgH
OTtDHtBzs0xjjoEkh2c50jU7gkHWU/ccSWfgEUDkPB9JwuWU/qNSJ1wbQ0ruX4Y+LRnWSS1a8XLA
Y6blzxB3ONpcQgFYB55MICf1Ce09jppH0sAFemh+YfM6bmrb1VLMZ8ggK/u07VxabQYYG7nuwPEQ
zTvAtLAfyjmSm3tBoIMB/tUo8daODzehzMjWsZDudvWp15L9J4eXNso2wqpnW9wEELaybg1x3UK7
z2WqNK5JTn5NEuErPS9xqz+pYYoZDnWYoJOKQPRRYbk1bf4t8T/J9aqvIGkYjPGOKjCSSTWy93Fs
jPELU5iiZgIKg583u84dUdJGWLtNOl1yfvOnKrJUwVEvzSjbU/IWaEN8sPWeEhDniwxIdTpFgOyz
rhgeICsueDIlvkxZByGYysH4ffx4KvnUk1FC3rm5IO7wDZrG2XvwUZxIdgndq4yGhtaWY0zu2vtt
NWnlLTgR1J5FbkMHhV4ZAQ44GIhxTgb2YalM1aqIfp+JThVU8GsRvM0Is06xXADGSpKnswMX6Kkg
HOCpAersV/QcRivVK41a4FKFDFM406S26PuzhAIrToOzpD9+21RfZ8pjvgLP1BWowQimeCD0yBhN
bVscjwMLN2EPNnOBckwwx9lNlFukU1921LmKxc0oPlSFLh9igRJIBJCOHc6LaLmISDpek/zdtTFN
7Jwsdm0jWMJ36z1yFGqB65bZnLzRhp55liKJ/GWlfTjOlFSZDTYSKZ/g7PFwa7QIDIAvvwKqcUzN
iqMDbc7Myv1Z6ksk2f8sp6abUVmB4/yd5PEFY4coc4JdAx1Cmxwm+RPXQMKRPkguKCcRqH57IHmN
MJ5zlPrerstzAh8MfgepxfXy8ROHU9ZkD6ATFiRk16U++XJ2Mg9X4YzP8kAKkT+Nab/11VM0NtDE
nozbnOeapEu68rEDFNXDC260UFb2TO0e9dGLKVbDXhlpBOUHNHbfRfVdDSTo+CBW8e4wCDHztjNS
rasj72Ne3FEXwA0YUBz4c2uWi+DxFkNNIpKEfslbri61UHB/4UvkFwew78fS7CPPvjoqYFfn15+Q
31XhNOCa6ho2+vGfocnI7+5OqVtgpXr4bE+U9b7oKmou+F4WbckXkOV8o5xJdjBrLf2EQbbj10LX
/OBwvlI9ikijzsEQojjz08IIBU8NSRc5Jt6KgxkTW05qy8vY3fjEWK9T080Aj3LLpZJHvPxoFPAO
swRNrDEczrhd+CkVJL3ts3hO5E46IWc60aAl5svzM3czlZYSNcl6td8Fzirw1g7az44jbSizVlA6
FBWe4lZCC/i2JRkrySdk4aVbYO3FOpz+MMe8wWwM2w9nOB1lxww8MT1U2pfo5ljW0fchCJ4wtfZm
4+ilDHqo5/ZNEZuZwVjIRniexUIdf0w4R0kt0OXRxpueLDTUiHjHJtAdTxCWjuLaDmwAEo7zRW+U
c7IoMZzwwWMFFS5cQ618H+BnlufwZs01A1S2fbePlOWlFmBRPwl+CFYoxvdz3uqnZk/gZQ4HNB/A
+rZNhE+J22AYXlOL27sT4NLtt7TFHdMMbkQyRrCXEGQGQngHuS5K/cwP6ZYCoBMYihnidIfyMdjE
pmDXSZFRagHFsWaAkSq2O8uFey4D8xHZ7dyXn/TiEZkMcq9i9ygkWmlmFodRlGOT/Z5KhmcTVU+K
RyoLu6VV9FFz+a/aLa6stz6EX5JFjMUt+kftJYIz3Cjl9mz3ciMZYijGlkQCyIKV161v6jPOAjhk
O8piMMzusT0urcG3KKCPMSEeNhmX8YltfSTc42AmQmZ4CWRSlzXYeRu0FDE6aagmXkTPCClHggL0
g9UTr7/wNg2TLazJJGGoINJhhCyujKIVeFwU2vvHDxOhRjzzvfnMHveO6Tr7MS7BLDGV5ZpZeLjQ
bMUkWGlhdRI40MVUn8UjX/PfmV+6veTmizhdrjsgXKlKzIbcjtZa4oxxLIJFHVQdyz7E1CNzzMBF
GeTBR1U8cUR0Vf46kLAN4aoZbF8Raxcno2SfYIBax0Wecrpy6fqv4AtwgG+uCoFU6pXaUE9VwYxi
E8YrrDQfVRtCk6JTMEBbpj+lyuBWk4GfciJfQRehmkgxV/bhlc2qAV1jkoglqkX1KeGtkbRiFLS+
vSb4rMPb8S64RkAKwKMfeiyMiHm8RYNqy52hbkBc4HhPTQ5C8X/dvafpU3MxvxPNgQagiUqIB8gZ
tm4oZoMAsivZI7oYOEUGI/IW0izBOPPmZN2Ik1Db4ym8S6Hy4BeDdUZxfMHxuxaqU/LTEqlqwXgO
bfPezTJgtcMick9mqRfXFltJoWrPFVctgEYjNkGXj8hgSyYQFk8mEp1a5gS0cJXqNjFU0dneVGeE
XAM9Fm4H161vCK1pvWCFJEL11LAQ0RWkd0ws2VzK8x8hH9IN0zpVO0TigsiCt74djpyVIObF3rP1
U3z2aiowQDZpO+6pvspl1e8u71XwcYDFxjM7nKcfaKWQaF5rOHVGdGk8Hxc4IrUh8BrOhNSsTA5K
ue0ERlYb8LNbXWIUF/rH/zeE+EG1wXO1an0u12uwD6TxkYaMxoYv/TrG/FYXBPwMBXkKVJlXejZH
loym6Bzk5lvEvaRq/RrMRUK9mwAVXyzs2TbMzAWZ5uziLn66lAvhFwwQZYTsQOxqtn8AhxIaYk3H
gE0TeFcVpgGqd+SCxSGR7dMFOWW762spgSPyTVu9IEvshrX9OMfknRj/YG/pXAW7jC9a4AraQ/d1
E/8gRv8X04+UELXTTeEENedsJ+t4Pq9j4C94iCxH4wQ/Av8VR6n8LY/VuxCvYghTKqkNAWJuY4A5
5GkuEju5dbpCpz5OWfyGsBf6CWajh/waml0agfLC/nE/WY8Zkm0dG6+Ml783lFX3uSiZUSFC+onj
jLnXaWsr1E6vPtFpWFPS2zjZdqXW3ITm4a8/wmd2lQgxFPi/0LxcpPxTTYPKygvNCd67B26Y1hoA
xP2cG+jVBq5DdbHn4TJwYPCcWTYmxAvSKXjPGJHi59LdVW/r3WWVkMz6QhONvW/7pcBZbpJZ3Iiy
YGqQRoTgadF0/ZjsbrhBLFG3ri4ynfJffFSqLUXYdi9Q9e40GHz913LM4ESX/1WT63DBFD5xmErt
0Zq7oDzabPUQbsV4XGiou2+P5PkvsMa5WRtrJWh0GUirIHYYR+BDOKXfQ3YF9en/rJS1CcZOQpX5
QnCcJnxMRN8/WYTf8eMneQvFiU2dRWLmPLKcXTJV8hVkPqATOlCl24K4XGDRjMkwQlrPkhulDW/Y
09odrNXK1JQvpPDIZ1pztf+8ivGYGM2OiJbzAY4wQ2DblhP4pNE9sCyCNESc8qQoN9g/JneEVeEN
mapdNdmcPP0+C900+wCS7Zlebw33hFUnYBzKxPYMs9C2jCbuiFcPxCkKbFBR/iU1Qu8F4V2aramI
aJjyxo+TY53U5Oh7c2Mveqm90ljduKDUODz00KpscpJ/yzKozst+JWSE0NDIQQUZTG+MN/ojpbx7
7XEd2rq0Tzb9OR4WGxR3mK+FvoQk9uy39gJZIwGPGd6+lBH76f+meRqacE1UnSpKuj4eZHlpGttM
GVAjI05REjafjl/VBLpBzR2v7wLgnnEieh5x5WiZ2TWy9+VKxSJ6NL9PaNbm1eXxRkqYwA9fwCzV
JUHo1GDhY7D9VnHaGOIttuAtfp/wr3z3QToPWmdnsHCd4ApWpWMVOvK6qmh/ExVbMjLvb55d/R1Q
NSvBmRchGdYg4FIZzb7MpYwbTPn9wxN/2zrFRuBy+iiu+3IENUvx0MWHEswNtphXz43/uPZsfwxE
tccKki+Oa7skalnGBOZ5DKkTG6Hn/7pMVaFvmJ8aEnu+efw5idunTOhHh3G9cEF2hYVaCFCfoTKo
JCh/3fMsqYQR6L374zX50khe4S9ZCMPXbUVcrb1VFSIYkYwU3K80TFZskE2yPUca57EAv61ZEgvz
fxOb8QxE6dDTyx6bxcLybfjSXf3yUFWX9Szvl1ScQgTh5/gb85gxKyGxnCBANjA0IuAS7f56DvWG
Oa2SGoR+1SGq+882W8DwLXtEE6Dkg5EcVr4A3okWxcsvFFUR2fIFkkkoAobK5uguHO6RZdtmBDG2
e46+QY9lnHfO7PPDo0YTQc/Ok8QzY3tbKSlQ3EcjcgT+YN8baDiPmKuOmTWL2UOo5LqXZ5Hq5378
K8G5VRjBz/buDteIk8e/LLUqdDdtBj7uQbFw5zeQlWNx4F+PV5Q6T87b1yj534hDN+lTXewdbrDf
1hXf2T2AxI1rYA08oFvhEceHhLFw7urb3XdXVDBwAwu3F6xw2AgB3UdgqWgeOH4/BztOZevSV+te
c8AegZf971otM9k/qzI8IEN3iCXaLUiLWbBo5+Xcy6YzU8agmoLJac5VBn5Pdnfj81F1ztA0dcf/
EGTwC7c86zVn7aTNhoJReykh3RMh34qW8StBX8b0ttR1W5nxffwcC2rLNH9RFLS/28lYDbdt2Clw
9fumigN3RU1I/pGYHh6qvSz9YJXX8SrEzG1JQf9gXW/B5dX2+ZpOTzVEoPuHe45wx8Q7aZygEPi7
BIAB6jSJ/ANthnKZj/iEjMVqSmEki3fC+6IWe569mvA/96cIcJ460Hs/r4EVz1ArOBETizjSb2l5
IRCqCY238iyazIePyak8FWDNbuCb2HcHrULhJSYyi9bHqI1r6Cw7uzRJUfZQtfAXYljivm2P+dsC
t0uqs5K48qToP9Yb//fG8dDjR5tfHjHZlxet94jH6xSOcSURJKyo9wXcq656MfrF8O4hcBaoUW4c
o9AccqBpaSsqD7Z4/vKunTJFUsveMyJeIdoGsCikGvjVWnu1wzoIPs9mR2BLUR9y3ek9JOR1c+tQ
p2cYSaW7mIyoMYzBnE4vE6KTNa/nNAeLZsEwKdo6YdJ1KfrwRcaRXe5AToh1hJPaocZFnq3Z7hHg
HDCaXDRm4UKDQAxVpB0Wwg2XhPf8lCb2qMBV3wDjGmvm3xODxXxUUmhkRaHnlrrib1FJtsEmGOaR
7anU3VpRT88IYRc2Oz2gQtqOzzMGUK1oDJYwLDQl7QPiCM4z1YNxjShLBdKokClUaV7L0qI+I1yg
EUJj9bEDJLt7l3ulNc+YMIRSXIWiJhZe/1WvyYZ91TsLqDHkvEXqFxIpwXV/VY/Vd7Mlpxbh9S2F
TQN+SowdNFrSMFV32seR2iwUNxFaGnPDoPEHwTSGyiYGH+Q4a63r0yZ5/jlRz72qAyer4cvSHiGv
fcQL7IObR51F5cbTPUaKbueKub+YQpzO9C8pX5oW0zUwifN1Iwk7Cs6f0oKkUb98oh0yHEaf1egR
KImy8lWn3wopK7DHTqOvvcQuEmqtt5AXzXsY9ZRGflXh5f85FripI2PMjFmBvg9nuZC6cigw0XLn
IiDEHZY2a3EvEzYh3PnLRVGTF4sbPXoE0LlHIE/ANFK3bwwax1mUeNDL6WQDIJIO+5HHMjG0PfXn
iIKu8tMaSbcWu8J3/B7oosPhmzJmxEI3ZgxMTWZv8IV7lh+LpH/j9hrd1y4JQCF8/8MCi18IHzB6
x8WvwSF3Ucgp3o4q6bF/hNPpQt/IUKDPuo16G0DvD9HEKydwIy6CnHAw7P6wTDVSOJAyi6CEwgYi
eP2TLIZLMQStFv6MvjwJ8w/WAvk7VOSrTrU1eMdhdfALI/SbpRerkh7IzAHj1c6ed2Kn9FHu44mI
iWCHwxVFHIdezwGlplNGQZ4LNUFItER0FC/SxccnHjAyPsoOeUT18Ma2oZhxDV8iu+kzgswdx5KV
5vDAG+ENQkywRqvmXXHLDBZa1rfCeFi3H9S6rgCbwfhQGunn+AIuR+vH/u+bNZTTQqg5jGnZsrFS
p844JYtVht9D4ejR4ucYic6obM9Dz1Ekoyy6Tx1qV4jaV0/TNVPUgCnrWTMRyCPXqC5Yowhkc2Lk
b1lsAYh2fiJbeAuDAUgDc0zbYPbCMGmUY+HnWsJMa+AvBCRVd1P3Sfko13Yklr9fXay7UK/pUMbN
OHzocMRw4s2YYq1DguTHCWA91Thvrrn946I/WrHhGiM3yqO8z5+XStGwnrRBh3xKLfMDXXpgw/ZH
MQq9E+SUryarRX+RbJ7DKtqt+pNpnw8bejRH2Wu2Eimdx+yDT/6a0io9FUTclU30PTjmN3uOxEpX
fouWFbYXQensJy3qIh6Z43RmDTOxr4Lqreo04oPtHtnxYbRdNlBAxomXkYkYt+NpzQeyus2A3Ris
RyibZzirH84sQ71fDdl2OJKdFBBrZO+qjhcUPYDWhGIfHZPcuQowJTb27krBDPb2ZRXeql94rue8
xXYaUfaNh/yeEx7ajn4sTUuq6S1DmfhZE/mJjn6bXTtktWN6lvqynMPmnlixODGqAmWerw4jwEbw
8a8kXz5ZB0oTWJVIHM28INRJJBMuou+PAeYInckd+++/zhY2VbogFaVvOhbeyBLoz4VXrGrC9XsX
wcmrTEon+JhU6BKpO1rwN2dLwKgzia7iljYQtp/SNhKxa4K+YpCqq26e5cKxG53m5l3EeONBVSQs
wrq4ncfSdEpGpa9HllZYzfXxJXQTXXqftpnateVIcpPdwSa/ERcktOzYRfsHOwXyK+S4oEyrh1ZR
B2nF2eHZCE4xlqr/IKZkveRnfGtsvrQ+CCCXNyFneY32CZDME6FOzNu82V7sYj0rxepexbnB/PRU
Ft6ALu6cCga28YgqX6cGvN2nr+vjfvs0mLadB7NcokPU7iMI5Fz1k9kTWnehTbKT2TWruZjRqy29
k8nC7RXOJracA6zCO6oiSb/tK6p98PIY3bgy/Ude7W6Q7anvLQ565lulfIT/fH4be1AW/7VwnFQ+
Vl0Eh3iLSZunlg+vSogqmf6HEB/KAbArA+Hpb0CgHAOBgoWd1bFFW2duJzYoaU/0a51+42pfTNqz
mXb7GpnzJn6mJ0u0rcVK/mClSSy4oGIfEZumYzZJdWWSs/eQfptN5URDAIRUwT2EibYfiL7OxGQJ
z+Sx5WwgWIesPT3DzZU8OHCmrdKN1RGLzyCDANECRoq9kVd5jAEmD0NtX8usqt01AiiHl0p+sIWu
3NtBK9rVaRPTZk7/j41TnGBhXlJU56tfWLiqC1VFIOLfJkQ3V3v+fYnlT7Uh//yamHkGMfZuZO5T
SqmdzDEWegKyYrp62yQ+X261UvPHqJ5ZbOJVvfs1GS8/UE1NBCH5bF063F4CbmE9Nnqlp3kg7Dsv
wjtnzD1JYiFWHcLJ51ZFikgNaStkkRo5TunQ7mt/YQlZ1zdneN/gYD34D4fMl3OivnhRyW7LZLfC
ENwuQQxr5hrTfBEh5xNlkPnYqe8gHZD1TWG44iFqszKIIjMpec8/iWpzEPUZQ5gbA0A6OmMViqT7
k/2oqs/UBwQbys0eYUQaWrC8C71XRKow1vteseOYbo1GnqqJygck9RLVKLUByS0b6lY/0VOjhH9D
W/m3XUmA7OmZsgRmxOGCGo5pKP3F52xzinx0qVXITlX7TYloNRbsUYblrBymwFsKJ+QsNoPVzZmI
06W7UvKVW7FJI0aFhwEz7V5jNanbd0Y6luVzKSoJzNF5Wcqq/L7V/mC4ISoAiHH/O/mQ0/Jds3In
nHqLfNA9XsGg+5m56uv1zyKOQDFdf6At+BFnjApN7tlwVCmWMVczLQj77Auwx0MZ0XjqJwWRRSqI
s59TAz6lzFMSqHvRO75t/G/8trzOPZQyicRodxYdVdPDVtGtHq2juGKb0PycqEgOD8dgzD6m/h/r
pCW+BJBxvXqSyFHiu236zQKua6fdkGW/EtmxOiRtkayE9DqRVaHmhe9kUN+lxEzfug6cdjOQA3lL
51/hanwbjjDL/1xf3UrbMDx/CPzKBpibuqnIR+xw16WiGSirVm2eaHB0wQx1hlsw3YH+1ZQyW4Wo
qVx63otrQ3B1uIawPVwERtkTsIUR+0PZS/LKhFGial4NCE5P+o7BYkuRQmMiwfbGPCSvHg2uxmUK
3qDRR2K57mQLdtkojrTU55s/YiPMu3IOqepvDHjDCh7uBn++U5P9G7eyiUutbuNGvHqWlikXxgbq
WRVHtZhShPbI8U5BEdG3tzfkIU05zteCqwpaSPdB6ATk8rLhMiM10Ng4J5A3mjpG2rt6LHG3fG4F
vOMsmPho9TSu7W0FZ6j1VitvM6ar+KoeuRkXFYkV9vbQYFYsFRLTmKqBsRY8eMABjb2TWjd1ku2e
A/oem/jAQct7nJ57ntf12JAfqbylJ60AbxaK9KCSE+1k0wIbhu35e47j27AMC2Qgv/3Xp/z+9S33
E11MHhaYaPrCPv8moAJPbnC6SZnR8d0Zs3Ufa4JbnCvbXWrUjmDy1t71XOoaEGCs6RDv6FiDO6sq
J5QLNYHKkcBSvislMnSWY1soHZRTuTUwsDlbosODV8XzXzj3fBXlIMvc1oyfJySUtfVNOouwpqwL
FHmqQBrPRBfIUxcPfrudC6s2H/FvsYPqLO7RidcogPUqR3+rQ3ZWmph6l4LRBTcdt5b7yi11jFEZ
zWbnCOsv+47IHk4Nh4XI+ZTDlr5/CzB5y7ZpzWr2lsk+rYLIty/SEzfaZX0o8erJc3ubA4f4sZod
TSQgh4GjaYsVYR830DFPgW/oAaXtlb0OH9mdDy2ZIYoKnJMeWndIpwVLTA2LP9HYPY0bsPfVZsTX
BiRx09SxcshQ08eV+0i1zgetUBd9BSQBf1ltGpP+ArmNbyy9OkmYq+0r4a42uNc5Msydyt++FXqo
egje7s5pEvf6G9DiSJbxOWyKD1BtOqPTtBlsQHloBlqOFCRgjxKjrb+URFAJv1xzEvADl7zJYVQ5
RJyh5lcVH0HSO+bhXwDXetLRnP1rs9GsB5bt5JerkK76wdGFSxcP8+wADCCpyJIKTXh/P+3iBo9C
+ofeBeTlY/LH/SfxsH6xomfUU0McTBcw8G705sQVi2UdVPc4oJctPaBWy7qYGoJCv9IcfdOzIhJj
Pj4PeJ4q97gNyQ7SWVGdkWIzw6xmfcstsMwoCTHEWmmjIZwZksKTGO42duF0qJAnT4Xy0dQCGX34
rSbudcKKoQzZlE2chFVy2gkFld14Flughu60RqQ0OLibEk2GxsXN9oubXS9SrCWU0AikZzE8VHv7
LoyhYB9B76g8c4Hpozc3hOyzyQxl4wPAccYUXVEC4ISH7VetGf0gmp439+CP4BmsIONGCl9rYTMs
oFefvyZw4warteu6IlnF15bPWUO/5N5UAX1TNj+bAZIh50RXQFp2fNMG4rLawGh459t5PkRxvtBr
8tz9dsHgDVaeZjYJzSGTXIuJId4sS0c4xfe11iopWir19xFzCc+cnp6eKxi5ltoIu1f2Io/vQbgE
qHY/TIvBtxo1pJTGfqSZargVOm86OXgnYz7gi6+iFY2+fFwZDWFbEXfIEX/zZTx9oHMGL7BpPaUV
uwgJw3xpqrtgZ52TJdqI7N0+6cRj5Tcbx1HS7l0reViQU3lbg0odS9nc6/ZKVvWiOKUYvh6L/0UW
m7+9vjZvoe25LJ9DZv7A9MNI1QMka4YoEnyxvXfBhcWWrBgpNg6hBInDo74va7ZtP45VjFI6fvrx
59ZhDzHMe2FzyYEWBJLGycvaW7ZJYVCrsWljNy/CQUwXQW5zRDeLuvgve6OxSuWzXZbd6bSWxUkk
8ax6Ue7weP3fquG6ynQKl5xtlMzHDork4+Y73/3oaA4H9/3VSp6XFLqrw8QJaTRmTMeLXPFUhDZm
knHpzSWKP5SDRUqErUiLNGYQbPeAQOcwCxi77qcrEnrQcVvD/cWQqw4cunUzFGqmYcZs6WTBO1Xy
dOX13/iGsRdk8tUmrFJSHYJTF+a/W/wHbM7rru88IOYrXNUDHqjx49gRUjPKZ2UaVkhE3YToHgHw
KK2QqqKgToG/5s2BVOk+c8rBtzQudPKzEMUyNlrcbmOQMyxw/yUZX2Mdc+Pd1fawRKDcYsmocmsP
2z94h94l4DKgrOVN9jZaYgMhfxr8jWU10dAgI0F3pm5Fp9JI/MH1lMlFGvnK8EBiXJNOtGoq7voL
WTwH1exnIF8/L9ZmmM3Uv/ecLZu9PYorwuPSs/lwf+HD6B2qJxZZOO2QZilFWmK1/pA2IBVYP5RY
HUGzYpYy9rN8cEI1JNG7oC9rL1g9sRslnFmRiZWfm1sOhNGJtPOm4zHjIXA/RX6iOzCsh++GwgDu
N1Dcls8hUV7qTjH5zfOvcrGgQa5M0XqxwOgYUzEMjeImD/PgEsCrhbKU9bUyWKoCsmb6ZfvCWjv4
+9j+OUofOfvVnN41oK6itAhJrPEslSmgJjopwSsWxq0jPA3qiGVh051QbDfbBU3FVf2SWprKOG/N
pjwv7fo45aDT+LATWx4d/ItSG3aTCfplON7JFB53tyT3pA1xSbGn5PUceMItRCCIrFrV7moqT9La
AoIi1DDQEmOE7MdkIrvivuNzvxHo7czCA0dMfrQTZaow3xiU5Y6thuOGFLF6ZXpZafm2eOti5NZe
1hWP3wepxZtNdBnURu74fIcvFFlxe31gahqFqKH/3kR+pv3bGZRInmvPd3sNYWUPrl9k4ZSLDR3y
tIfMBOJu+f53NDvLNzEL9jEoNAI8FW7RfvxhqKzJPJsYdgVJRDh8sLqDG3nTZ8YdIwNq+8pErXpg
tShfF6jN1fTeSIDjsEbAC2yo9i51m6dYjyZaU4AGSISllrJXfiYhVjq+gUj930WLvoXToXIQOGPS
bmA/TF2qBen/iBjc76ByQQtzIyi4RgrkjvCu3PUOx72ZhbOM5rPy/RbuBHhKUzpUPrMR9XJVmYBK
cTafT/NABLk5M3F8QXmibe2/Y4fPB4xXSyZFkp7y9YA9H7o35cL5J4F8P9zFb0fHdhe+hmlWQPQz
J/TYzdN1i9MF2pwFaZ/K9FIWn8wl9HopaBaBWKB41B+Ael2dW3kT8BS0UTQUYpC8XWL+Grcquymc
UMwyLL6PS5k6zuiUdJVwcu2P+acbDs1MjB2vh3IFNQkVJT4PXA0YXCq6Rq++rJkTOapviOK5unLW
D+boZZjVwZVAx4QCosW81p2b3xYJwleczL3xZ2+zYKE8PS7catXhHAsJxGbev++92HW7E9X4SLPY
Tb7Mzt1xNswrQUIhZ1Pz4dHAH9949WAg4DE2ATMW9sCUvZDOLIky2a0EkrdIuwfh0yz94XK9bkmI
KIATefpaXTO5hddvrE2Htl3iFUZyw6cU7avxU7mLUg/IRt6Ey4AfQtzvFd/I1i+vyrS0x9fA9TBm
SPv8KnKpruAKt+w9U+8qarYXCVacfxg6r/YSCT8JmaBK7q2cyxOg1mmTYWP/H0+j1wefeoON3nW6
cLfYiR8gMxmlVXwFcQ1mFHXOrTKHgCM+Sivxq76TnTMX0CJEep+fjtBgIiiZ5oLVUzXhIGAWRtCc
9hhlgccROpQRbQsbT0A1TYKrkr5guhq/MQJtMkxgSBbu0y3rtOBazTjq0IzbqjD5iFYzArPrgPgs
qduG8NkeKjkeKiynadXW+p/kDFx+fErgddE65uiSodDkVkHqYY8+tfRdFJJHXAR8I9pIUwj9YWLe
zhzqrp+x6Gn8+UJBHK3d5UWa7IIEQ56AtwVAEdvugz4N6z1ftGZjthsEhTeIILDUMq4AndVO+cOJ
9Vjturz27AR+pzIAfc5vJcyJBUaQ1R/S+sWJZU8Sp/V09M59dIr1pl0dUfK2fobWd8Wks4NypYwL
X5g9Ke2unLMWyqZ1NDBMV+H/Chaf6uzm5mr1mbN5SNd0zpmE/xwAisLQ5yTUvg9gKF1MJ3sD4+u+
6Csg7DeVqnp/RTToqMuNHdDaP1itfOTL/ZRXh40ga9rRghi2XJ3nQIqDvAOZZ20S85QJUgd/RR5h
gn2ss21KRFZWeCi5Qo85pZ7E9LS/Vvpy2AMNvBvdaYzJhUjJauZEHP7eqndRqwA2xxLIQvZG9PWi
lrsby3gJnkmb1p6d3ugnjAsIOBNej1IUjpfx36SP8TPmw7uSgAzmv94mETk6IewenjERDVhsAx1C
WExpaEgimQl3WuSNqnLYHulgeXf4n9cbJMduBMagDIKd5n9EB05/Kcy35cS0XS/Nf2yHpF4lZGTe
uELlA1aKmLhDi9Bb0EQLtHBQsjuVmBUGSFp4XUL589Uz5RaToRjhaZh7XaFPA8Tg5FKA4o2Q/pSA
+8Mu+LlA1X+2WIKdV9VEM3Kj+duGpJqOH+schPRrb/LV2FqIiiF5Qcw3F8V9GzjMjFAd/q0zlC5F
w0DIoXKISNHCxpeCI0jZCY1Qs6KajWvyXVKlQ2aGAX88lbVu3O0fdSPChM64WKR7qO6HFeLEQGHq
eHS/kyxrjhVWvuFYAyNFAdTQd4TcL1igG38q0S5b7c5+zwtqZanVoGpeTaedbfqf0fzmXbFcyIRO
qTKMKTWs2P1ABHFP+yhViF8TnaDyHHdw5fYoUNbq2URyk59HGrM9jPPzcxC9BqKbj6XH4U8vD3Vc
lFMVPEECKwNNnDtabmC7OXBt8Za3uVHPhqXzA7qpCaukWzwZnwY3D2Gmx1qx16mzjp0ZwAxX4Epw
Lsj9GADumIdC6uqmgl7xmf3O/q/nVlz4EvkncBCQ9yubW06EpNL45FFmxGT+vElGdXD9kym1CliC
aoY2BBMVu/Ue31lUsw9HNFRbFJhpXCienL2LeoP5GNVpe9xV3isMDZPdQDMuD7q5yzv61PsJLFG1
O7B1M8fUtziJjzZarluRXWGbH+20oX3y/xN/R1+nEXSqmKbM+o+Gz4i9q6fsZ16UfvczDmbGPr5k
P5HRw7wHyqKbhx7gLGTBU7PV12mpDX6tw4rOda5TRqmUA+HpnzGHOpXKQufNhMTos2dzFyNwNPXx
XQZbCkrNQd8gANXRmpOLpSo84AC+K0GUCIvwRvZW/ARfSHawIvSYI08gjlTVPZKR82+h7mDd9Q9O
vNUNDdh/nf4fPMSZ9vyK8kc65CezhaefG+6+8PhxOFJuYo4AU2p39F1sKvzXb9/H9Zny0YX5w1MA
0W4XTOgfUgNw/pDFfyL4LoX8F76mj+icnyW0+trZKmtHQC6G+sAzRIppOnmn75RW18ebh4XE5fWc
olchnJONEhguZmz7sahjygKyZ43Rsg5rzVE1TCyIjnMjy26HG9VMF97egs5gytILWt/g/8fKzaGe
Ryb90FxqwbSiZCvpYYGbF4l4QnUZg2UuegiUKgCsCw0vsgAxPoI3lbGuDeMBhTJRAYs96EQq6C2P
QD6pkl5L+UOmm1O0TzMSsffT0vbdZ4MHF4FvJwLQR5sefAibJQFE3+qC4+JlAxfm5hT+isZEbluY
wT8TYrhs9JxvLEVmDDcI9EEjb/J+r8KO2ZdHH58uN9oG2VJ4k45UfFLyLNojB9d05SttannKvS0w
xrRG1dfOIF/pdwO9RPvd5f9dL62lA8XJqZSudztD8Ohhq74qnM7fq7ZrOSPT/4D6Wc7/h+uiwzu9
1bWzAY8Ac2LUHToidMzcW5n+zr8c36bk3qrKChuR2kheCAGmAr+vPiSQoiZrKkktti3l1KJ7EKnr
KLaS4pDk38Duf1pB1aG3ZDtAcGNGxwToC9FruaKr096T8909OwOfC7Sdfi69LqOpk0XGPNOkILEI
E1o+tp0e4YUGL6tdpgFysT0EaboD/jevMWaNdvoOkXPAY7wRU+Wl8N2NNAgm7k7712W8S/Egv5Y/
6Zauj1hGDrPq55qN1Tzey/ZYLH6SacdY4oOHWzEXAiPNrrf6rE4SYqT3IAZLqehBTcH2VKVoLBcm
pIGSEVyIS5BQV6ztt/mL+RjhHcCem5L5I55taCKmQvKkF5Kfz9QrSYJnijaUOzZ5Ts7VBGHEcgAM
Ke84M33F+FNIhQY2taIwqSAX6MCvzAazohHbENjGxKjLzFh3r/kpbJANiI4NukgJ44ta8PzmBc+a
8cfrzZI3VOCeRymSW9y3yEVEJcPFhHEdDO20wppkWU1R3yMlF5uqwmrJe3JX4E4FPBh++eURS8D6
G11l0WlQj4zhJ4vcxgYVoSgTamKvHNoqAWkOc9XZAcH4lFYAma7IzmlzcFmlzNnP+rzf0F4aVrW+
0ToBOH617mPtKixaODdWovKUGDDwJY/8kbTIiUIgX1js2oOYojPWQboCWibEyJ4z+PBe2HyOYnd+
joZ7Gx5qonF/LMCvwi3U1LJthhGFZwNRYvb+4hbsRVFf8XU7uRm+Zz7RL2CT6JgtL7UJySNpjcZk
HvNpUd2ZmJOZ/78A5J92TEpRhW6YrUyQhjobMR1Reo2GCna+gMh+3KXS4PzO2sDu+nCErtZK0fzO
/sqhxzEoJrMsX3/Pccu0MolbVKlB9zAeqrkmC7ckXzfK/xDHSCBcLfn29b2cjl7dRIOq+MF6MsrG
5RPRU1RORTCpk7TWDcNeM9LpeBO1qrBXRJM9CouNZETj5sKgq+S8C3tguCKvBu0L9zXDRGObyfGt
lV9OjGazmYJeuON88uB8JDaneWVmraUN0l4AmAe7ugzbmobiXZpJF7ZjK7i1ZvDKf1y+RXdTCbt3
QzOeQZSHi5cCLl/mL+9f0z8/FV3OJtKMqiHiyESluNFKKmI/bfZOk7RxFiNpP1PTb1BS4KVPIYn5
bT9gSttXjWuH4vV4kEyIIbtw+XYAHUKZkctMvMkr9+BBePOGcNBzHskHycQWqNy3FRgISVhfUiUu
5XsZ3ejkFvluSds4ZOa7oh08XzU9Ht2GUPIl14dioLfQieACmjn2u6GNoQhw7k5A8fZXnT3S4pAG
23hCFDwqm+6sY4rMgoSCEIGp2LrQCXMh/R2gFbz30UjAqmS2XJLbC5sfyUm1R02bWMAg3W7Y6Gwk
9LZVOwVXo0aB2rUePYS3JBqS1HUXBu4RgKYO6YCg4JjdCwTcA2phqtl7MArlgMYG4AsZ9BGJIxze
A65vAUKY9JXCm9Wbg4ExbhlAp3l0wCShQBxl/vOL2R7KuUez5DRaQfJeeu8QJS8hk5hINi0Spepz
KDWX+Cpnn8Yy0ZXUUDnAJ21h8gi0knQvQyeCQkDt5c5RhS+A0kX17NlZFNm1t0qUcqxIOaoIzw49
UFsvxhdDn/HO/EtihWqsLIOg0/NbC68Ex0xAS2MOL5XlXoNydBniRmgl3fU+aoeUoAENsG9yeTs4
UOUcSy3Kf+1flABP+Dixyo2dSGpEwR9/kE6USNhNdCBkfxn3gaJODBeYYlijjRrmS/wMMzhhh8G+
rOXEMs85jail9VwWqFRvVK1oYs+4KD6QFvXdgExtXoHG90QZHl61AklSkShg6PGvCX1JUx7/eV1/
FfSRmFn1ijUt0dG6OoCk7Z0Vq93glUo52hFiE5VqrVzevaYzgVTWH0fMe93iXMac2CTUzM0W3fj3
WPwALgIK/PCNJ1xPhRCY191V48UfUTczsCAUZkK1glLxxMcjuSY00DDPhtF7bRLCrjce16a8NDKM
a3pMHnpIh6YMdezeMhmBEERuIIpz4s3H9EJh2R0VDjIuSTAP5poFfZ4jnF5RAWtxlL+6XkwedRGO
jAA3pBVG/2ymqQYx5LfbWmToegmzaVKBeTE9hcoIOJyoH5Z8/UB2XHAvJP9vtDYkvUIU+XQqMZ80
RYlMNQkrpj/MYaUEZYGLloD0fpUYD7gj//y1RmNoKMXZGNRATU9+rnZJ2EuuBrqYVLukugItj6l3
3u8CJ0bpML7wgX7y2/gwJTNlAV42boiENrJBZL5tsNkSAdhFvHEavyZlQYTOq8CdkU9gDNz1tRTW
1mcahGRMfzQ8Gk89wCPKjMTW5HY6jTXoqem8LnIFEzHSKHrlIyRFKT8uNnNQZQia0zqfYwwYFYnH
Y8sKEx4fdv36XEJtefwJzJKbReQF2kxihQu4EEaZ+kSAOyUHd8zUMOghQddO6rNmcitZ2LRZ86wH
1iNXOxMWRmvadSXnnkCiUvmhn2UpRfyHaoyLO5eObtwAFLn3Oak9vI9wRtxiGfKSRfeUNK3eBZ/+
Mtf8xXXUWlBWo/BxPD7s3W6mzteQaJK1rj/dCUJQqMaxQRRjV110FOOXANTrTr3modj5TRV+C98N
kUhbBEbMK54R3KLlxKHXLusriLH6KvfJi4SJMGFJQNttKmb/cSUdg8N2r9UzO42sRhUIeaHywdTX
VypGQAKmwV+TqdAJpkoJ6PEpn4wasyTl74LDKe4djAIQJWWy/QwDRHKZ2YduOHle+ihDvuAaFNxr
ltrhig3rFgUhi9TL8mTbmcl3g1UkT92h70bfzR1wQ5cUAMBqeVtnco7ddyH2lpIcsoYZoxDZJ/dC
53Nd0n6wRIhFbRzWNeK9Y+jbZBBtGgmeUdYt7Zxb+quGw6aWtsLEkVSKNDZAilTr0H1sMz9YFOZF
qdUw7YRQRzR9LZWA1k3HsqpjjOWI5e6FAid82ZsU0pp5Dv8YOhUxSYICi7jDoYodcfCzIrFyg+kR
+FyhCCyB4gP8sVedWT7MsPkeW472+FSLyAmDACdA3Nvr0rwdKhjA8R3h1K80j8liBksFwOc8RZK9
/Ybc5Vs975KlkXkmVsCpT4balwGT9vZ/r0HiVDK65iKnYbGlpUsK15hS7r4NLjQwRtFVkkMS1T40
vRQk8B0MY9Bs1M4QdipSpnftey+RboPHJwyzlWz1+DsoT784YxF4nh5dvzm6aVLEiGjk7C5WAyTF
n4xszkoXbbBIFTdPCqw/oBqeGn1UtHGH7LEKtSIQyPnukG5lq9pIMIqMIZ99iJSNFE1FMQVKVnVS
Bx1uDMnylN5KeMP/kisXhYDWKXApUpQUgxHJ2nGjX9LQS1/2oaI3Xig2+H1AxAP0uivWvuSjSFAX
UObWk9yrYD2kYX4piKOFmvq3iz8Vp7+PJDtSo+7OI5mynx/nacplJpx9/FaeDHHNHqOvlgtRrdvG
uMzUhajSz854khDwqFLuOm7qFsKcGjA/IURJDTr2dpsFt8OzY8hMasZgh4q4MeKxpJOxvLBkQIXW
Xj9w405rmivzSBvTyn6mzRSJo8GSyqm5AnaS3eyJhwcL8fmS5/uvuImYHtmDsV1Ij8f7VSXuw3zr
1JX8YmdBKKfgq0yp7olCvShgL61bC6xj3veljRCZ9bsqP6XAdVCKz0zs8GWkKqKCAxx0tONdxcOO
zWjiRI13gxmjhPYas1VNAA9Nc4WhDkv1R4g92CaKF2BBo510GWkqaNP2Zql4IBJHiGTkKXyAF/l7
yMMNqqjy10E6v1oCYXUM7irR62D9uPT1m23xpdMZgZaVjXfg8n2tpfkZQQgONSLoPzWSygvep3Ai
yo3rU+4eYz0vgBD/59/avCmaTottJGdeReU7cMERf3M7FQ9TT74UWx5RthpLdmlXYkl2asCZ5P/8
iNx7d5NekGyRRW760nDbZg2OJ5IPTcgfl2gpwR1u7fB5W5TvGlP/z17nrrd7fHc7vRxlykEdwa+G
IVjvH/MR/zMSoQrWxkReZz3gB+u5jsRAADbDFWVAxfU6/+QRlUiGDhqx9D3Xh/3zX7DeyEkcvc8v
bn1uHTtXhpApkHBMYM6OWxWBC6VrB/Dq6imr/3NeWTUoCXw306xIIXr8xoBTZ7/I/SmdWBJjp2AO
p7ClnSC5sT+MScgHkFeVzGgh71wn6zS+AKHNDdBJS6c4hSmMUVft2vDcToyRCHBMeJDS3hnIfFBl
5f5JSEZeW7XcZstEx6VRsN8d+hFNUWwip4ZGS67vjC2Lg9xR9SvAmk7stOHXNKTRlKvGG0SK7bMO
Twer4KDdwtQZ0QYZW9tvfm98YfIUP2UrbBGgrawMuxyAxLZjO657GBIFQW4193pAYBA+7025a6Bs
s3gG3rcPYeMxHGRT/0xAydHDBx4Ok3Or/SVdWFGQzFmzLNUM9aXkboEW5DXN7URhvaw4TCiTyulg
gf/ixH4pdnpRHNn0cDIAwCyyqfodUK8SBqLRBbhqhDYONkMQAcIMtxBsEudATwQTcecxS9+Ndmb9
qd0NaJ1kXR5By0IoqpTI9b6EhaK5TQBEx+PLNax+8MOpShSlbtTZN5rJCfJ2WiHFhNkzt8EygJ3d
YTj0hA/FXPmpEVh++vvmeALj1Pk6UPVhqbBdv+qEGTx09u28ZmbktlGV4D1ScZKVxNTI49E4tKBw
jD6buA4a07/Qen+AiAgmWkFi5t1DqkVYCSJ/n+JXNQ56PRn+QjOa+j4JDRyLZY2FPQ+JrbymIHGp
KBcTkkmIiZIFcuGPtiRJ2IBwt98DdDHbRJKNO6rP2Jz83MU3hAVM6fvEgKOkxzhvlOqFjV+e8mTK
M/RaPrMK8PDOO+oO5spP9h+nlIHeokDuMsx3h6317NrL2AE9DQYY8JxRXItgK2cErUbYu3v4Zm3+
mmAJPRFX6fseKG4be92aP1+grTaK0waAq6Wh+9pje40ougyQyBwlbCZAIVHN5M+wUK8DEqN15mV9
fIhHuHp5lQwC3DEbZnwGcoQmdWoejie6dgieuQODvzBLJBGRACWxRQPO9YnD2Q/h9c+SJZ2fLQE/
KP3Z/jqqtztVR5mriWwiZ9jszbxTIw2NX43h3dTqBvoBG57Nli3mpTocIjQ1cIF776VdmksIFy2b
EUDasdCCkpKLG8VeeOacVTPdkRd4DH4KUJc/GeTFZCTs/rnd5qYSV1Tt7QRxTWOLDz9OPAz/Tli0
QRdTAglIJkh0RCNZr9Wyv3/WznqVp4cufvcH6Wwy76DdsQcEsSVKMY84ZlQq+KjuxTu9c4fl4fJC
KqtaHn06rP1XOTU4s6xbUvlNOJfaBt3zPG2TZ/rdx6518Mggo1ruhoU09Nh+/iQkD7mBuZVtIRL7
XmtL4taaOPAS3ef88YvYFl3ttdfy8KCbSPWs6I3jp4Xrka1vcODutBa9ZH06RTh5WQs5d/PD/ETp
0IdhV/v+w3JTmyzkhEBCnZKdaOuMQKv+8xer6La9MgHm4GAVZXdWiZpPLNpMrhOGL+fQjOSOqTtm
d9KZJsWX/12qD0py+0RTt3L9amUER/ZvSNlKiuSzNiAd+U3u8qQmBg0YZVm+ptBC4p79a7NN1n9O
jp1394ZJrlAfbqPwHYcMsKeBjiNNL/Xzrc6UGXnXlNc/VdfK3AhQH2XFiXa/8/zA/6mCOWIDXYe/
L/zqnY4/qml/Aohd+wDoTl7nTSocGecOVGSnjfyUzJe3JElQki2X8gceVfk5IKSxKMG/nR79VREC
JKxRS9AWhX2zmNN+/QDosfQMjk/4t8zkVEPF2HRA+kZDFRAj0rJolTKBcu0q1gRs7ofw/mtgqLO9
OknWrfVQYcN24hk1nQ4QPWeCUKCNtc6+Dvl1XlcdHks38cEnuhXJWEQyTFiwh3asLy3iwW9Z7gyA
lz1FQXiZXOWYNk2wMhkIuBVsKA5nucsgDaCupUtouz8WLgY0e/Lh2W13Eln0Jbah6UqxXn8b6m1U
DuFJrB0j4wcFppHIsNMlGqV+qtWgdwbaYNP2ih4mejNuftTb5F5wpb9YBw5997kZHurTn/xZ7A/W
+EmOV7xZiXqSciarIUuiioKEl1q3v7JlFDgzgkwEkSHyVxJ2PTU4nj9affwtpCbuaf2RHgmxzOxu
UHuING+Q32WdQqBNTopG7ps1MxLfsB0T9wEcH7H2SP1KIpJNEXC4CjRuSX03G4ojvcIh0Ioisxzf
bzYl2oZzv8QFcj+cUpz+RxmvgIkKDvZMAXW4YBRwUGk75SKauWhzXgmj9nmZaEKW9xKKcn6ppjqU
apAkyCmJ/mqlg/jjW5jX5FWD2xHgQHLzQXOCJKIoxvDDtBld8Dj/LP2GNeauDO3I8YJOmckg4WvX
U5DKuIr3SzC5/UaF8bscIxkD2vxMW34GCEiD10B8JPkK034dpbN2DKGHn0hTrhRNoTiZTe/Xg0eX
MTO0XL2VChWhWdgnce/ZnObxPnTs0X1Y+xx5AFvCw3xYoGqEfXzsfztUDCtdtHNtnX9HSxw6wsRj
0PKo9yKZU58ECAedXDW2Nb6Nqm/GPYl+A4ipdmwO8hzhn0MMsRuTpQWz7i2uJHdTHOSN6e8hTh2B
h2kBwkg9HTuO5kmvF6Ww1jLLouz6nJ26y9QGbOWxuLlj9xHXfKkkVU2fgGNRq00YQmkaIcB0h3nH
zLxpH7UNf6Z4cNMa8gMxURZ2FRsNTcbscldytWi1mH/oCMb6XCz3Lymf4aIwQknYLgEbvJsevqM6
ftp9vEErMi/Qcq1dvst/uQhC4RmkPJPyDvaxd/A4wieHL/tq483YfyTBk7oiahcJGl6K0+NwTpe4
HWDdfbI/usO4GqD8rw7/Irew+v3KqDpFwXmjrATqWT0e0ZeUbsSafI+EHl+NWqOpDauvi4KB0XZ0
o+gEI2O6P3wrBc4hntvzWcfVPfhkb+q0XK9uNgMx1OQLZlWaeFllQX4qE86kFIdnBNJ/Yf1WByYf
brAEyDxphuyZHTHMeTw7jsWCS1LfQoB5epdtKVDA2IMdnwTU3UaGl4+B2YpXA+FOAV5jpwJajHIc
jXEspDWedQex0V1qamLmzszcQ5/u73Z3vPMyxo1vDfOKmaev2cueVTrqDMspWaAiho4AW+aiNqO9
rFHJ4lA0m7kmYF3/ki3iUrz8JxAtjwwghnSVytGkQdaIu8Efo4EFEG9T/Mzjo8yzJZF/zy2rDiOE
l3uVMTGAHlv530gKQfG1Wvg0y16oaJ2GK2JPnYW8Ekn+I1OVYo85NaOHCrDOaORUJK4m9ED5sziT
GmmdcZjDFSR14TEAFuX1oSDfyp/bVE/XW13oKdCkUy3zW2awzdsNkasH8qRgTA0E+K7etLfNSfYl
u/TB09xpEb+NH098BghyVimhNkbS1SMwnhhfufUG6xOZn/S99K0l/pDuFzDmcDTK3dyJ+TI895jY
oAIQ8Nl6EfV2Hpg/y88QSgPuLSPFdPpAAYslwHwLe2muLggFfiSFxGNV/quY6cGpaD4suJ4QR4Pr
JZZtyDrWUw69gWOcsYgEVa3axmr3Fza0I8p+W+GEO+hq+DbdPYsw22V1yKEKS5qjhxhBL1zmSa1w
mRZKsbreO9ZwXqM4Gin2VgEF5YfZeElYKzkoSHHaFXJHhCSSY3oib8aQa1xlxrCvnUm1cnHz/k0A
vc+5qRRHLvkLYuTEjoGFVCFKdO0ZpOo/bftJBquHudVzYI2EhCfJaNw324p7od7LR+HbcU2NlEVB
WmuTDsaORbtOpyUSgvC2lCJR8QmNCbFOWzzorPT489Q58AEzPrMGgmvIIy7Aa3oPETtZfhRhw6l3
XLg6k567BLlvzSQniC1qN3iqXGO2aiE3b4wwNGgqk8mQ0/F+OXE17oq5eN33R9d2tPZ4H/T42zTF
+bSAT3KRUzugECo2epUU6Ninhuj0mV2ZTZGZhMwst3L5pjuJ5/ybBdvqWzBSKza1A9k1kopl7lKN
ytG9gvxAjRLr6rKt/9yMSdW/+GJ7JbraF0DU8OH0pfTvEhHxcQIOpqNLeAnSI7Rluxuv+resQFPD
vcR6ye7UsWK+g+GhC0ZjQibTcPsoPJqH4zjb4TZTHoiVVsw6zVv+3MkU9/CuBm77J+5N5GL/LIMU
aozJHR7XiOwrQfzuDbgUyQs1nmKWqn26KtPrZYxcUfdygmptCcrs+vEyfGVALL7f0jx7X9lX2Sd9
vuqoF0DvOYHXUWMlGcMUkQakiTjDez2yGmbaG8ok+HMeFVAWLkl4/ombj/pOpL/SqP2K8/uQKap0
e+gfNSbAD/CuomxNQm1Q/LWXtLNUjpzMdNrv2ffqMxiQeIxjlxCMpPbVmTZQe+Ab9Z00do90PK31
g/xbWtibdpi0aPj1XHMTMxxm9iVmeh3AEVYzDRm1Vicd7+lymCFmnxoVN7cdd/HfeKkLezDYA3mY
VyJ1aZ1Y7/G7pG/n3dDTEp8xrCBHImI0qvzK7Gy7b/Ym8NksQZy7kDkmsWUhR9kJEUl62ECiyq6B
kmYcxC5bGKIcN2+uHCB3RMTxuPqFui5OpbzIT8J1hnZQ3UWXauNuagOs0dkXqoOZvD4O8NmvemQb
qErxnjbM8LsmgHbVhQbT5VQJDEo4788io9EUL3SLvz6ojU2vVCNrCQz61UmGJ4Awg9yG6NkiLput
pfpdAWQe4cXb7u4m7xq9E41SA/p++nplgBWjl+jtzminc2G2tQNMcJKGiG0iqQ/ZpOxpcJP9t6tn
/iA2VBXyn/BmXHkmNAAUZGr4z/3wEQOMhIBUoZJEX7RNS3CffOHhvnlVXOZ7ex40u6pSIBB1zgDv
QDsh2AwvSxDQgDVxAUuaiwUWTJTj71uQNZ+2FcY97VtgZTBHzH3WC5b4oUdDqzEBTnJtBAQs/My7
u1XyX7KEQCy5eGAbYLHVjtXVqDIVQg/0frRXUnJfKgxSHqFEE36q++eUItleT/tckj/zmwks+7wv
J0EqYTqObI9a+DUK7w/yN/LOq2DpoynMsQjxhhbHpNKfo8cyYBF0By4Xe0MDCEhnTDFkDOEB1H3Y
CqkMMaXBjjyZAxrBgCOoWTV5CeQHev8j4xM/n8XoLlx6uvaIAn7M0krPTQaS8hgu1IBNbbjImHiS
1lT3U9tVMCtFKWy8MJQql4WwAHjz5WynDGK0Vzll1OJDinJWOdkivi/zlyogapdBg+MJHF0ya8VQ
OVQoJ8ZNrxAXEo+AS2gpQmXBDn5wqbITMo1ySN62feB4bKUDCOdgtfB4YL9NOnsNL1TDlitwL2LW
TX57gAIJlwg4x+vLwK5GOCeZEBw/1kn2iiKrTzexBoRuVGOSvZqVzI/vLgyIA+SipVpM9ZjjfoWS
dG24C0SWwX1TD44DQUqI+Tb4Y8o5QFP58eQGmCKQxrsgWZ59eoX+ChWUPPfGvP3j64vFLCiHt1Fw
NiRDPFSnD7yJCb/vhMeqFHHLxsy52u09qt+gPWJI32wJzvuYOMXx+beIRMMzZx1GtQJ0LZahwJui
wnwDtlryiWc7+vRiCV4TDsIRd5eeaMte8M2OwWe52jL6GS1M54OFgZRzMBtr8KDIiNHmRYNoCQfh
i2Vr1hGLqw0t6VrOxefhrxp+hQA5z8xIV95ZumLqGqwEOG0h1AzXmuBlwbDr+jy0CpT2KAuQf9M2
f/20e0B2mtYOuGrzwmGCvfBGMfsRK2y25B+2urOXzEq3ae5A65YKV401tfFMN6KxKe7EsRydFI7F
52mqLBcG4zxS6HIwGF3sluzf2BB+E9I5E6/sHVPuR2poKMXcJzqpMlAP3sGNHsL7vUd3nmVapKSY
ae1HP2nJNXJ4bCxx6vAanVtwDJv1ZAi6ELVhW48Gbv4kC30o3rbhu7fNRWxVpNBkRiyvSXncfnwX
y8n8WIDvQdb2NsuvApnvAxdIlLAW6mbWmXueEfZOJrfXdVohQK8r69NCtOu8Aguomut4LQN+nex4
P5TkmVaYIF+vmtp1uWl2+lPrz/7SLfgd0nI7mztUYY78fq6uqQWLEimKANVLFP91eAtRMXBTYgJv
xW1UKVITJUW6QH0M0PtRLjBDlVeDmh6mcMdTrNbQgqk+HOLVTGcgbQpaz6XzcnN4cXcASfulLtds
bN/ESMLCmnc2YzYfpBJx9gufmEjK2vuCSCR0IGa45xY/fny4gK3dgvHQ6Bp0iyMbMIN0f+xnUeYK
WuCAR+aoRZghROCHYiIgAVbzMFVxXx+Ik6JCMq++/6VPUSu92BQxCuKPRVnA4H0Irs8K0D5qeGfy
+Kh8B7iAPbayS++ZU7/ElIcVdXMnrqfD2dO5FA09TwvXo+FRokOBzykuEhGvHs7OgEVSwOvAClVc
P+iaEYYyax+YqpQ2W9z2OXtYKZvCamCgXpWs9yJ7XHkOpqPi2reAZNLWL0l88JB2y4wRvd/Pt7CC
lySE7JO7qwCl3Cvug5F++j4R/HV+SGrMtH4mmpk+NcEX46Ur+SrbpPrXo0FOmcTwt7I+T0PijnxT
1IElnJietQtATCVdBIy7vv14e6mRYURSzHdE+iWjCMLi2/wN77xx9l+AKRy4tuGVrcQGpZAKY+Sl
++jjJeop5mZUYP7J3CNIfZFK2YKU8GwIGDWiiz6L0Grh9OtaR2JRaq4oohThufyguNkWAwDbXwYT
3vOqumeh29tcT4902Up1Gdz5RusQZufeqJrvcavVtma7Hp5Q2TYOvqTCXXPBXDf90Fypqsb5XxgQ
cPUqYlKLLKKrtMbgjsDM0VBVIy/7Dn7jJ3UrBAecMLnOS/9CnSirxYlesx4mjMW0wGx92tb4k3B5
GURGlVug3/D6gjKpbZ3hIYOabMVeDTN+sd7dtfdSYaUAOWUCnwf24EwNJTqYDmyCfkDKLK808a0o
AhCxOzjM1zNTaaV3VhZml/npiJM9HQ2dfQ9OcwIebultRqwV19m95BakFseHoz1EU8VrRBoCFyVG
cMu1SQfKiwgWaVIBsjeDwKFXYUWp986kJLDV0UQHw2+CnXEu8ctoN+DERJ2OqIne3enjM0IGIqEJ
oNOcQsGeD2T3p9a8jm+99JI9EUVLT2oivU1TL0f2XueCHG4oCrrwiedJ16n2GOTTishk+AdTTRhd
7iBM8cDbdNKcXf9oyU0Ex5zaHrDSatfYzx+Uagd2PYh8GlqhHruwwWRh2PoHAnFbOU9AG8QJEanU
osN1mkwMD2vfX+P/DTK4gjd4Etq8wC5sIL/vSQtIKCDy7EQCNIDUK0a99zbI7n94pSNm13Zsf52m
1REpQLqg5WvkHSxpIgls108S2FSB/IMRwE3ajHjJoiSFRKYmvGtw816+PnRcIB+LPAkfCwcjxbWc
q2sSjYfgnar0oeRJC720uQARYBxZWa+46Sibrd3zlyH5+hiLrz0LrGQIGfhKEvmIYRR/GptLcxai
NYXm7dcGmgJpOBaYY/aSY2aggREImZZDTrtMgdWnSfV+yNM4qauGFEV1GSmTS8CHQ5QxKBlz2UX0
2zIoO7Ihv+GCRqIVa/j7V8g/mZI2HiGWkJb1YDXU6q+wDvWSDukuHdWOrUKpEAZVeEHqm0dVEal4
2Lqcgvlm4BxxOHfbsgFnO+iVY93+dN/+L63ZiSiIFNZyUWhBk6MHigbduKlRV1dUv9vDTx4S0YYA
3+uZj0XqGIxuSD9ZGMlTpAJvHmQ5K+pFKp07/LhuwBIhvWwgt6+/ayQTMezEno3gW9TXOOBRW80L
c40XsHs8YmJfeGbVWhY7tcI/BqQUTHqa0cVsKuQcW8YbxuQyv4QHnd7lh3XTk14lWmb0fufRDcxQ
H3lzKjdql2hiitT0ZPCZ1EsXmAKl39xvsiS9mELwTqBKgGbudwZxsWjiimwX7Q5kFFYIUctLtWOg
rb1B91Fj2bZl77Gq8IHPgUUmmuLE0Muus4Gq4hqrjvtd5OALgaUsAfjnNkS3mSMdccskAwg4+WG4
VIIupFOUMW98Q8+xmcvyRU5PYsVBmfI/7ZKcH8fR0tGV4jlDDodCvkBTwFcoWsko9xifv8pZn5LN
fPNMh/aNjvUB4ujiBc1skrjDjuqjl4J1hX3OtoeT/vAuuYmBq6GerySnxbaFOI355RFRCvybcuUu
NQK3MWKLrPA6D/UKBtWfVI9ekzArqGkpjq+0hoSx1WlOQTS1mKccwjB+A4IAICdW/e/nNjfAxHzj
ql0JTLyreTsBZr3zLJyUx10Y4vYYe6Jt1/UQvU3hH2w8BbhRCPFOWyQag6STQGTZno6F80HQLaik
HHRK2ui0hP9XggvHs1hO1HdPtI5O4Nug3K3q1iFpEmkKgmlklcbg9TGZ7ikBRH3DWLHOk8YFvO5u
dHqsSg9dVmvIgi550DRFZ7ya1DwQODxIXx779glOVv74fr2FyeDyRjp10ufhkfjkqCtVxfCudG7s
bz3nybqAFVA3IJa+YJWEodHIjwSGWFMCTkZTaXjUWgVFDzBxWDUtAp3kl9RdHpOJwshphlaqsd33
PyUY+045jJaHgEddgqH+BuHXLvi2IjSqizuTb6KuCNdfOpPv1Mx+VvaCj+Yn4eaM43YYrk42pcuV
x8t0LG5pTlM1aIhkFewytkR51Pq0dBZs0w2TQBoNY+q5e2ldlWoclzH26DtlVVScOWzmN4AjpPEq
NPwTvkftANTpvMWdXyroo/y6P48bCsRTk12pDjBIJY2m+OOdaWRX7pLBO9zjsPHiJ4bF2D+ewCQJ
y9sNil4ygOzEa3ZWDrXHF4t7rnYPBUOE5arVTv0PfPGnxMuttq7ffuQl4AkxyigfCYotFlWUnwwu
n2aWP+VCZUrcgLnHP0pOsBfe2bMYNnWE30nhGTH+VXTwFFGeQ/+ziW29pxto+bJ9vPN4Ek0ZKJXZ
+AKKIGXKTvwOod9As/973a/hcWB5rBX00HXauliwgP2hK8XfOrC4XO178g/kdfLVzdYdnZ2K9+BM
+W3/EpxCohPwE6W73QSb2PCR6vC2qL1+2MADlPfdOi0OXgrK7+rHxR52qHhTtYKErvFru2agQIgZ
lOE67wEqgUnpu9XMhpQ4fk+OoOaY6FNlqXti44vNpvNOknVoAIwFrHL/vGmDPGiU4WMQBQAdD8gF
fMIhZjiItOtByiI2S4IoajegyyMWZuz66/Si7dSuLOXraQuPsH3+aodfjkwNyvS9ewD7Pk9fs2z7
U7xgHZo/yfHseYeWifBqyoIAto5vqCfuFsRtSefE6LBTwCiGBIp1Ipguen/VfDIHHV00H+tZF+gm
QuT1aWipGws5jaowxTOvmSEjM0ZqpPutkeV8s3jBOvYZn0NoGuJYXoKx9KWNKEepwmbIFI+XlEop
Hmlto542v9eEkfZajx7Sx68RKKc/Hs6KIRAC+T/NuYcjuiMwi1h187dM3rSFVJfZw9uBIjcyqYWj
ESw6sob5VH+3NFixLnoF+c4EKa8vf16GHuaNI7CLtKJqTA9HKVqw0BVddQ5sY3fcLBzyYS98N/ly
k/QZX3TseLM9aAh8ouKkUr4CAFOSwyB3+jFr0U2x23ETyD/dJSadm0UBn0g+Yzadpas=
`protect end_protected
