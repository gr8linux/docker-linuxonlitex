//********************************************************************
//
// <File>     : const.vh
// <Author>   : GOWIN
// <Function> : Constant
// <Version>  : 1.1
//
//********************************************************************


`ifdef CONST_VH
`else
`define CONST_VH


// Module name
`define getname(oriName,tmodule_name) \~oriName.tmodule_name


// Const variables definitions
`define	AHBDEC_ADDR_MSB             31
`define	AHB_SLAVE_OFFSET_UNIT       19
`define	AHBDEC_DATA_WIDTH           32
`define AHBDEC_DATA_MSB             (`AHBDEC_DATA_WIDTH - 1)
`define AHBDEC_ADDR_DECODE_WIDTH    32
`define	AHBDEC_ADDR_DECODE_MSB      (`AHBDEC_ADDR_DECODE_WIDTH - 1)

`define	AHB_SLAVE_0_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_1_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_2_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_3_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_4_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_5_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_6_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_7_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_8_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_9_OFFSET_LSB      (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_10_OFFSET_LSB     (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_11_OFFSET_LSB     (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_12_OFFSET_LSB     (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_13_OFFSET_LSB     (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_14_OFFSET_LSB     (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)
`define	AHB_SLAVE_15_OFFSET_LSB     (`AHB_SLAVE_OFFSET_UNIT + `AHB_SLAVE_ADDR_SIZE)

`define AHB_SLAVE_0_OFFSET          `AHB_BUS_BASE_ADDR
`define AHB_SLAVE_1_OFFSET          `AHB_BUS_BASE_ADDR + (1<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_2_OFFSET          `AHB_BUS_BASE_ADDR + (2<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_3_OFFSET          `AHB_BUS_BASE_ADDR + (3<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_4_OFFSET          `AHB_BUS_BASE_ADDR + (4<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_5_OFFSET          `AHB_BUS_BASE_ADDR + (5<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_6_OFFSET          `AHB_BUS_BASE_ADDR + (6<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_7_OFFSET          `AHB_BUS_BASE_ADDR + (7<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_8_OFFSET          `AHB_BUS_BASE_ADDR + (8<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_9_OFFSET          `AHB_BUS_BASE_ADDR + (9<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_10_OFFSET         `AHB_BUS_BASE_ADDR + (10<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_11_OFFSET         `AHB_BUS_BASE_ADDR + (11<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_12_OFFSET         `AHB_BUS_BASE_ADDR + (12<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_13_OFFSET         `AHB_BUS_BASE_ADDR + (13<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_14_OFFSET         `AHB_BUS_BASE_ADDR + (14<<`AHB_SLAVE_0_OFFSET_LSB)
`define AHB_SLAVE_15_OFFSET         `AHB_BUS_BASE_ADDR + (15<<`AHB_SLAVE_0_OFFSET_LSB)


`endif  /* CONST_VH */