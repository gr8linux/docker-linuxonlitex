`define module_name JESD204B_Top
