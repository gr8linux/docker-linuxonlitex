`ifndef STATIC_MACRO_VH
`define STATIC_MACRO_VH

//`define getname(oriName,tmodule_name) \~oriName.tmodule_name    

`endif
