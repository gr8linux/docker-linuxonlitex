`define TX_AND_RX_EN
`define JESD_TX 1
`define JESD_RX 1
`define LANE 2
`define BUFFER_SIZE 1024
`define RPAT_EN 0
`define JSPAT_EN  0
`define INIT_SYSMODE 0
`define INIT_SCAMEBLE 0
`define INIT_F 3
`define INIT_K 31
`define INIT_REINIT_MODE 0
`define FIX_EN 0
`define FIX_SCAM 0
`define FIX_F 0
`define MODE 1
`define CFG_CLK 10000000
