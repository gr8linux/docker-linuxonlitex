
`ifdef ADVSPI_CONST_VH
`else
`define ADVSPI_CONST_VH

`define ADVSPI_PRODUCT_ID		32'h02002044


`ifdef ADVSPI_MEM_SUPPORT
	`define ADVSPIBUS_EXIST
`elsif ADVSPI_REG 
	`define ADVSPIBUS_EXIST
`endif

`ifdef ADVSPI_SPI_ADDR_WIDTH_24
	`define ADVSPI_SPI_ADDR_WIDTH	24
`else
	`define ADVSPI_SPI_ADDR_WIDTH	32
`endif
`define ADVSPI_SPI_ADDR_MSB		(`ADVSPI_SPI_ADDR_WIDTH - 1)

`ifdef ADVSPI_ADDR_WIDTH_24
	`define ADVSPI_HADDR_WIDTH 24
`else
	`define ADVSPI_HADDR_WIDTH 32
`endif

`define ADVSPI_HMASTER_BIT 4

`define ADVSPI_HSPLIT_BIT (1<<`ADVSPI_HMASTER_BIT)

`ifdef ADVSPI_MEM_SUPPORT
	`define ADVSPI_MEM_SUPPORT
`elsif ADVSPI_EILM_MEM_SUPPORT
	`define ADVSPI_MEM_SUPPORT
`endif

`ifdef ADVSPI_QUADSPI_SUPPORT
	`define ADVSPI_QUADDUAL_SUPPORT
`elsif ADVSPI_DUALSPI_SUPPORT
	`define ADVSPI_QUADDUAL_SUPPORT
`endif

`define ADVSPI_TXFIFO_WIDTH 32
`define ADVSPI_RXFIFO_WIDTH 32

`ifdef ADVSPI_TXFIFO_DEPTH_16W
	`define ADVSPI_TXFPTR_BITS	5
	`define ADVSPI_TXFIFO_DEPTH_INF	2'h3
`elsif ADVSPI_TXFIFO_DEPTH_8W
	`define ADVSPI_TXFPTR_BITS	4
	`define ADVSPI_TXFIFO_DEPTH_INF	2'h2
`elsif ADVSPI_TXFIFO_DEPTH_4W
	`define ADVSPI_TXFPTR_BITS	3
	`define ADVSPI_TXFIFO_DEPTH_INF	2'h1
`else
	`define ADVSPI_TXFPTR_BITS	2
	`define ADVSPI_TXFIFO_DEPTH_INF	2'h0
`endif

`define ADVSPI_TXFIFO_DEPTH		(1 << (`ADVSPI_TXFPTR_BITS - 1))

`ifdef ADVSPI_RXFIFO_DEPTH_16W
	`define ADVSPI_RXFPTR_BITS	5
	`define ADVSPI_RXFIFO_DEPTH_INF	2'h3
`elsif ADVSPI_RXFIFO_DEPTH_8W
	`define ADVSPI_RXFPTR_BITS	4
	`define ADVSPI_RXFIFO_DEPTH_INF	2'h2
`elsif ADVSPI_RXFIFO_DEPTH_4W
	`define ADVSPI_RXFPTR_BITS	3
	`define ADVSPI_RXFIFO_DEPTH_INF	2'h1
`else
	`define ADVSPI_RXFPTR_BITS	2
	`define ADVSPI_RXFIFO_DEPTH_INF	2'h0
`endif

`define ADVSPI_RXFIFO_DEPTH		(1 << (`ADVSPI_RXFPTR_BITS - 1))

`endif
