`define module_name Uart_to_Bus_Top
