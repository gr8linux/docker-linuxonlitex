`pragma protect begin_protected
`pragma protect version="2.0"
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="GOWIN"
`pragma protect encrypt_agent_info="GOWIN Encrypt Version 2.0"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GOWIN",key_keyname="GWK2021-01",key_method="rsa"
`pragma protect key_block
egrG0DiLDmVP33C+e3XMbkoX/BSW56Hao6GntdYLFnlzQkRzk25hrjyt/E0zIF+6LInBWJG5aDtJ
sgtqKx9QOQuS4wojLDMXc84i1SliMeHyUX3efGGZOCQ4c3gnPy7/r416L+sr3kcqS3Pg/LiEP7O5
4kmZ9IDI9MkdtTv8sEIR63zORXIvxavkJVPzmYGC42tYmZpy/dXIPTOdaLq2kx9eZoPyk3B4xpku
F9t7+0LX9JTpXIbQrJYUA3u3F/M1KQC+ww95ZIRi0JQo8RtJ1w1iVIXOS+slfo0fd1WiZiJD3S6S
8zx0Oo9tIFB9OFmvYyB9VFCBw4LOzhozRHpUqw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=117504)
`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
vH23gc4Hv8XwDNbJTi8GjvxUBgqVGSV9DkOr4HADMWOU2wgqBFGccdSY1xnjkc3037ZM5To1Xe9H
JZnP8OSBNyySxCpVHXn66hha1Vi/fDCZt/FAdh2HCleAtLcUMoJUnhgxGcCCTj/TGdse5W/iegn5
6xjWSBybQg1kPCdEbETIlMwsPQUjkLI5C4b6Mfc1EqtNyV0MCcFmHnnctd3NWvcq7IK3dfEJwHit
OBLKV871/2NU3NV6HBgCv6A6YULDHRr84gYaF8JOV7Ja/hPq11ncdbMeo1F3caMQY9yf6lZHuKmW
iCzRtBXLM6h3qq4Ig2IDGh6sNriMjj/XIbf9w750z8T4keLR2hlTAFAa9lSu70t5mf3zhOfIAozx
o7Y+kCdei3Q0Vdq6QHDMhWz5D6YSM8SXP1WB24H9T7FWdgEeL0PVd9o1RQyqxq12Tl9a3TkoaNRW
NYFyXEZ8fQS4B3fr9/soxPMUd5CY9nfEa93k5BBbLTHJ/HO8795j2iHZMadKMybVOVlFarn/VdZA
xur1CzV+is7nKV9KqXnotgdfseouRX0A38/t1mUf/RkBkh3PjD+8HQ8UC85zNjvKVrpe2K1X5EpW
vvMRZv8KP0AA2P/Z3IFmghMCAPG43kjSVtoLK2r1RjEvSyncj689TLxEejg42Mg65IdJHg2hTOIt
iGfVREjBrawWOrX+ejVvwRt47wYi7TXukXGkWOxIlyXfP2qukVw/BGnHq9IgdH/HUnkEsXisgnYL
AUnMKX8SYsrptXPf3r4p3xVFO3p+1ffKooYkUOfBXKC37gIzWpCAuDCXNAzCQov+PMntHCnNOPdG
L7luqA2Kr6mc4E4fZjcWmmLwpyOxdFdtugVPzdwqpKBuWC5mI/Rlks9QXVE5tJHv0PGFIuSe9dy1
GLdcPk6BCgwc1DzvyV7T8zKRfb9HMAJgpBYEqPJjJs9TMIz5zvizpusRpCfvpkJ5mLRgKb30MJ4M
PNRVSFCPDyYwBml2wONcJ+pqMnzBzZ7EKCRIfppldZBH4NpG12mND/wWYI8Y/l9buMyo0hZ+wawK
PuM/UnJA+2qx6Il4NTsQ2316UMPFHXV2gV9Goky+sFoib7LwXmyZ25sgfEaQ9Vo43qQZNcCN/0Ve
BHW74vUjFxyBtqYYfjNlQJm9UPbpD31WtEGl/VKJ0RzvT8YyFvNyTTKkecq2y6tQ+i7Gr6dIHAno
SsnCdS5jPNhePCndZTF9a4MlvwMKdEZHRKUAyePVVAnxkL6bYx1vGI3HmgMFwV5vBtsMa0cQTypg
oHx0BxWfGe3KJRMPX8QlfsY8irBOPSV2wzXxk2M1HWuZuPN3rV06+/40YmGhZsSIPtq5d5n4Ew4y
EPXUHPwOx0LHiYr4VVexev8RfebRdQdnlL/rGEVhoEnGSQlF35YtT2H7g/ONDMo6++fx7zW7Xy8g
LgToKCI3Ey8QQHlqnNpAxFgY7j2OgRJQ3xcYCSBhFrMqherdQ8GYe30iNvp1L0+LPX2SqtcfS856
F2zKOJnJA8yXMmmVw1fOzx+oVu3utkAuQVVUprOt9cU0q5l0Vsc+eEZUKDck4dUK6Zeg6EFBoW94
aLvvEOiRwcWLXT1bGA/r4kH9kmNrtluHwFIpDjl3vJ8XUdne3kimdRNhFM1/+Z2YBr3699PwzyQL
IhHzXzV5WNWZSFBbN80voSjzTcmVewpABtlgr0/3dChalKkflNoWXpS2Ibs/qlmNZkr9suzuBQva
WJXHAJihzpvAsGZOPHPn2hUYHBdGJKlfOn3WAXO1nluN84hM4uHXbZOFpSx6Gtj67op6bDAo8j9L
gRUBKHZ60c7dSISy5tQxPLBs5WY6pc/2/ID/trTmBBkHdzDoreNkDdO+fcUNWKwf1qWMDbkgiGtu
mXzOiJmy+ygRLJEyWJA9Z1uXS+FvHJZTmYuY3FnkJkl67qEuTHgw5HnIKs4O4k1LQbwnuxYgDZQK
FIlVvsHIooSPWBie8NvWCg63m0EwfGqpBeHW4hLs+1Xu0HqbRI4eY2/1qttuPtiZRsc7j+ESvVBe
Vt7ylM75IiX9HQxtytfMmi7MtHkCMznNE+THJ7bRLuUQf1IBFhbAOIbmKQyJF28VFBQulOWXL+j+
ZGxrPtVRiGIHcbiQ8FLmCJUZyDoe16s/Ta3QVQYVuuy815h/JX0/l6/g8+jcoxeZKSgn1irrlBNP
7d92otvhPse7CXdNe+9jF2QBIQYGx4HXwAdSmTagJMsl+paKswitSKkBMxpafZfeXTdNBtDt0nOm
P3MD08W9DYUoGWd7j+xCgd9a11VcLBuV4w+lpH8uUvDBXAz9VrubRwwwThTrjUiKoP2YgxVRvF/F
jNHhpIVD1E2C3Pka9FbKtjrr28gSELr5lsvJb2s2Ba99DWnuNqSWQKsTqWHg7If2MIWAu0icOJ86
ZFp+466lKtUo/kS6hw0oOmczaXIpjQiiOYzBo3mDFU1bt0F1SFohUD5jaqEv4OVag36hBsjS2bwt
IWCfUAaBBqs3Z3bSIAwJi+Boa+WjusuOO14BJSyD3/zXsAZDhNRY6yGMDSsQzdt5dm759FK/IhJ9
6JxpspU8vKj25M/6O+KbjmDTJ40Tbz7Dc1K1B11mEmgQ+vWuLI7OHBXNM/N9linWBZlLrqMkKFDf
VoXXbyegKcPv+Y0kC9T/v8NRxMxMilDeDPnBlXyQdiDvFjDWPE53Fssvpr3F3pRqaotYmF5I1kQ8
z3E/6eRS+RuCKVs9o7bO/BCxB21fST6++XLHRyNebjkyPwOfMg4Eqc4DxHksN2zvbk69alLBbhZY
ZD3xOkRnScbdjTknwG01qOTX4ahCptYwvO9fNJfvyojvGGqe2A0uZ7E3Uqc6dYCxE2s4y0kx9/0A
6a85oZeOGoU+YXeTrLIjdFm8zjxDpPw/TCgSIcITBK6OJDre1sefmvzOdNR9kPPP9VmPMnWfB+GH
c/l8P6DBCOiQXEXFbvccmo9vNjPBF3I3C+3dxHUYCyoQ9TXVoB3OUgro+aQAUDWvd3m2zoSeGgu6
VGtiVcTo7PjHf3NQ1GxtIRf5Tn1qg08dQhOEaRoQdOin1ILFlmGI9aEwBRns/vZjtKtT6gRzAer+
QROmEOrXbVLtY5+ujEeRZRrcSnNavi4d7OvB+D5M5ecPJhV4cEJIX5Y49AWD1DLo5w4ixVA9C2Ez
064q/JnPmkGEyyv5hVMabsOVz+5SYp1qTspg2czRfHj9zdjcrcoShMEW8J+50CDjSROuLkJlETep
8w0P+BBXvf7bRvAgIfmI3KyPAjTkSTQzkIog+/5AlWFXbVBEP96/2V6FR94PlJNEF8vpth9RoK38
qehgUo+k519RvGG669RMboX+5xQaI08PVTgdwPnuynGU18tsnBuO/GCetQoxqGeAhfFelR+YfhV6
c5twzNgPHa3C4cndi07rzxZaUUyP17ZlARI9T7I/xHgqHN7ipMnAnB00TZ2fzlEgR7PIPayRDBtL
3zqXRb67AI0rwbJCLTXUDfaeRAHzJxUiswp6BC2qLQMhwj/XvSXgPJMz8eW4dsrKHfQf7FLOAICb
DWscicGYDNOyqgsyu3+ZSqpts5AOVqDJW9yrhXyN9IbyAA9yHbyWBBDY1WCphEqjFkA7San0Fv4H
sTzd/RP/iv8LNo/yl5ib4iaAbvxHDW88ED+LSZidGFccGb9za3WHD8Km0NMbSN0a+tz7KM52w1Xf
6NA17P7UUjLJje5AJzk06bkMP65gANmI0WvfFZqfyHgJLlq+c3AQIENwVlnow41p6o/s1kAsgD0V
rWe/QFAnAxF4Lrrhgp+oD/etd4ui/FX9T3S0Raz70KUbcK6W8B+p9urvb0n+CgstAAdRXoUnLWfd
Vs18nuZrMYMCpD4vA8Q8ZKGceC8JaidcIuvdtshyz6TUi6LqUlRudgKGZHow5iKWOjFcjCx/6NIb
CJA+9M1h3sn7dS6J7/MTZvDPu7hcGlrsUK7vO8YnVsz/jTLlE8eotroCPTKaJYI+kQXPPTaiMfmb
SLsNHByGFtM+4H9qZGuXTZ5zj+BxAuLa0JMlMiXT8tDMwTb2fZL37w0nFMAwL+l3/4OLLB/eqV8M
5JBgt2/sw7n8MrrTbdlYAh54aoSYc2T7b+UVTBwGk6Rm2E2oKEIw1lJD5f/MptSjo6aFhQfojSx3
KRJZj3PxhdH1XE/mVaoq/C/dMUST0NmZHR2japtoz41VToro1uvXYQRB4wKL/vWFS5RlkdDCXrcN
rJvQsu7VfHicjJCPmdGs0eA9rAHea0r9RN7yr7rwsPR5VT0CXChBjDutvlXEsQi/tXjtdTm7xU2S
uxjWr5kjmoRJDbF/bGi/QORIVfzsKh3bYkHalsyBNo7kCjZdKm/9iK5sefmas92e9LGiwxqSUmYy
jUDIMUE3UtWqggW6hyqrLYtlF66zOkm3NwRrvN12N56k7YyH8FC3NzvUAmY2gOqXAN5sclyvDifd
VMU0TPfEGSj79gtQYptbWaVD4i36nGDJB9h1kSV4cDUwvBfIjFwrxXvEv7Eoc4wZ7oXZi0nbEunx
WdjWngetccX/Lt5GvKjpA4eeYCy1UY99XC0H5eFmztvqhvOKcXqai2JcgmmdeyE44F8gANf9iavQ
shazwZgb67JXtMCFlIUKyCIa/5WcY7Ig5faqXHWQ9gsSlVKvRe2exeQ5ERope3PPjnBSDbf+YP/u
SckIjeGvxJDa0O5riS2BUB/j50xdDWFxZC7380Mo9C+2TekIwx0ny1G0B11X/27NL9+s+2Vw0Bao
ZdxaoPNUPj6WQI094DBdx/j8zMXwZGUZMDRQ9fUWh3zDcwW5mVM3gOpMkgi9VI5G2dJVbyLhW3eN
v3mfFW0yFIV73yVXh/drQ8aD/665ogv/FPvYh61X/xpE7IlL2vW9GO/OxCiia6jGTnLgS3orIS9d
+Li2LeeUakaTTrsux8sNLAqCBrzwws4X1FSPQCg7k/5BleWng4IIE65UPRo1FMilPL8tJtocSwgE
wHf4GFNivzS59m8jq8loanizhMbFaO31MOhiyu+yRxki1as2ZgbSMQeZg0S5Odb8ToElUUCR3jRo
uwzLZmBByE3X0zv+6+IrGwVNSniTydCeySvvW7u5rEMb06RL6GG1jOMTVipDIGDrcU3+u6AcNs6r
0epMQoRqlgRehOo8GnpOMTFuiaO3h7C2vJoOvQ1UVQsakN5s/N1c3bQWDYFZSIOzbA+4mghTopEw
1j/2WUVQHWmBx9JhY67CFbtgtGuRrAlTpZCcCLtNRmnJC0T3fiR8xwiqXWnyhvZFa9IvfZPCbtjE
ZwAAj5b5Q3zy5E3Fbsc8S2pGc6mkbQeWUiDK/0EDTKinWEFpJbbjthv9GjPn3agyBFsN9SEHl5cX
vBsWoPFI4nk+myRHNKyE9FxTkKNK5C4kYVkAorYoO215p7YRly0hN8wOzPEnCC7K3Z9LX8025NhV
6UzM17GBxjC8R1zg4cLdRcNTih0bSRRohP/AYCe1Rf/FcoSXhV5SktWRCa65bvXUNpWhSCqRlOBV
dG3R0arN1M5roWPxNW9v9q/HceCh2O8Di5OAMgfeeyn7wKLhUM+u3o4VqG7d3Ou81daPzB9utNzr
CPfb33OPBItWT1W1c4HCCJwOF4RB+au3jq+++gdJPSgkVswLFhs4VGPn5boXj1kQZZVRdFKM6zgL
XccDTHZFyIQYMLqkk5chaU0lpqQT3QgrRsy4sO3J5ZwW3gQgHhs9tbCB85ze5mxUBP/oCAzJlCKy
UemnQdt3st1mDbqj4B0hU1Bfqm+/kFtcV3mdn6DkJUtVJNPF7K5GeTrVCz5VWW/ZNbZADQuzX6vG
qltmTI8U1DS7MHY8iVIMM4t3M9gUrIKfwrrrTz19MArgwHgCHOrVyVFsmYEO6TIlNeiyv5fxLEZd
eNqrbTjgxNFZTl5uQ0wwEn9n879hhYO/EvObNx+d4iL5XmuAiI6MFvQPKyERkJ5WFBo736TD8L9q
msOobTkY2n8YwKpw6cyaKT/Wr5yVlV3mDZuyRDtY6u89p/4QqjyRGDUXXSatJ2mIkvlm2go+xhFQ
fNtCsVcGdqyEuijfX+e/5Um9yF6JT//BshZsNeEk2SO5QMJlkhsHWL6jV2+5UGTKJ/LE20YGqz6f
lrfenDFqXAG5SzRKkiFbXMZlvusfM8Wy40puGo1R2qzeglxL6XtjBqSowR5Z8NMrBC1ebTKgFU1F
cP1e5K1Bhi63eVyK8ufcgKCG4zrxegMNobGzEVm6HX636fUdVsLDu+3rLBh3tsX1S+6K/gauwOv3
EaXsioQRrhtR9Ywsam2eDKBOj3ogt7QXNFeJewfbke3AfH9RGqhDCI5pOUgP5y1feJSS9iDyQ/YQ
drNMYcWDKTRouyr2zap6wFiVcQMgm3A1wwFhWN2g7IoLL8qVPSA2Qp9j7QWg4AhB3GfaMrXwC6NN
86Ko1kmfJ291pJ9+pGgEdvp0oqYHL24F1pzDQfI7OL3H5nzGUxJsYozirZNHZWRf5bLG3wIzVTxj
NAhhDiy7gmLdG5L1rjb8dV9cMjAte+uS1yc0Dg62uLlMuI+XLOFAnpegDwjxAnuyl0EU01W2LuDc
g4s1CPmTzVvJciLHQepeFPeEbJgUJrValkOa7e30t1iorv4+OPhTnbXe2+qvcgGGKc50PiFl7/1z
x7P4uuyT0iDY1HctDKy1Q0QaKsIl1iNVtK30JotKKvpEc0sCL19D6WjK7N/OkrvSlEmqNL4+aJzt
KvQJvu+WhvZRh3/Ic+mI4XTYODVQFBXGHOzL9I9OH98MllIIE5RB197cxTlso+wXFXNgR7p720lu
T5I16dgTOsKLUYtKS/pI1X7MkxSh4sPHBnFMAjAvjfzBKh+kUt0/6CFl2wNUPUXn03e0mp5D1YUN
XYJybgncfikWzeZdHMlkSVEjbVospQ/7Y47L/zsYMwJXiMSFGBCP33M4nXLp5y8X8gOM02KhUSsy
uGsktPJx1aqJyiSZZc6W1lGJDMfY0vmGb5xIeIF6XHTPoc629CUPRVq98iIiGSUyRJt7BV7/dErQ
i2ksnuHjgmAwlUXDYERXnQaMJrWYdLhJqcv7lNNRgakcdbD9SqWxzxehiFoZPdewUag/SFsjEYU3
GB6GgtOMQ24YC0uXzXdwnNaUW/OBylg73ZpSc0JdZEpbF6vqG4by6MW2RxvxrkpPmQ90ggmG0I7b
C/vJr0gnaPrikZ1OM7zQCDqze6C23gEw+Pgw04SZUFAyaQ0vUEXcDYWbFAAKuOgEF5ZC1zIL51Lr
TRCP7d2Dln8cqgDLAWU4gSXpyuu4cNNx77zYVd15/lMS1ajFqrODI2zRKnqtAIllGyBNhLJ+u2Z3
qfpy5ZrfyLznBetWW2MqPz84gQxIviPnJ9DtnjuTjfRFS0TjvNx0bdGBFbJ/5Grsu4AmfzT8xwL/
xxIdF7Y0JUgNknXspkSSrLqZGr5CyJzQ1WFgszKbDMOOcoScaiNN9LUzVcizU5BA6wAMijdaNtFW
GBSfVfCOTKatideYzKTFmsTVEsG2WKnxSK/LL6ora9r9pSXKzxf738oH02IXDe00pL3zT3gd9i5e
gr3JvSYzdJYzCxsLuFkFg0OicQ+gqqy9ZaJe6dQv6w7mV83xgeA2CXrws19+3Fy2JoxlNiyz8ALv
1yIZlw+IKIzsaPSuH8vSM0KjfsO7StYIFZYGy8sQX1nFE1/wxXGvgTe8TpdV9+DbdSNXbLMHzHSQ
8J6iuQzoIYx3iAh3Phf9mA/ZNRZvtPAtSNrKPmsxsuciGiBt2ovZsPM7Xqy4ktfbAZ7sQ4e0USHs
FqARwq3fyXYlK/kMuhmLa9X9xs/jKm1RSOYnkcBYDx11aQIKFwWuTlrgg7+Roc6xA7+lFWoOBtLf
Y3wKYIZ+ylCzP5kFEoHr+/2FTWsRreLcvs36zA+0mywAp5jkOzzdf3LRwuV9q5eJGC+lGq6dmJsW
c+cm5cPLHZ8RmpmuPb2TEoO+UHhbK2PWrI7V8/9y3eobVR6gojVdPAgIqUXstnXAOVg6DFz/y4/w
5oWMLG5F5S2zT0svzuE1qKrmZxrAkGRfj1ac++1T8LNurZG/QmdUOZ0+gihhcuz/AArpUUv4ibyU
2gSx5NQfRQDApFT0Xpb5hjU61YJ8veCKR42N4y3Q/v2kHZLP6kmfryr+EMWljnWhaQ1I/9AaLcGY
iXaO/v6Q+LG17BDIuFcMnesb8FuBj4bvbIYZ2MGOq3e/htzrMPFG57jzDF69gLL+VKVSVMfH72Ks
kU+lM5ehx1U98LJ5CW0E48G0grYQWD7/RimAt7QrpF6fV6hgaUEzJzIKD1LzjaTk0A5NzSZiWNgR
bykWlrkxKIkCQs7Gjo3y5NhQ41dEUziv6A8/dqeoDI92G2UK2ryUfbGbyUegDOBG7lATtKRJZu5k
k+8308lAB7ixGRWiTnZ3E566vRCAJnsoImPIOTx8n/7OiVargTPrd/ZdhgWmCseODVsG+N+TEMTy
m/rtDaIZFsA2SdhgG6UAtPx4zwR/IqibLDnXdyOlk1etY9B0cSJUL92cE+zH2k+a/NVi4QyaUmOd
MnNZEXhMAkgZj2C5cUB7fVBrrRRfHkTokXd3egMxwUy0Rg7yf0CzLKa2Nncexq55CjL8I6Y7fDI4
zGVAhOVTYOwHslgSw9xtlfB5QI4C0J+A1HjDIm4fTIjt1FlS+8wsWjPLx7Em6Tm5PLQE7vGiDlP1
KlXFb46A9iT5KFUgJOT4Xx9OjpL1IClUez4kNsRCZGXXdBBEPtCw1kRyf9xzpO98AH0mFdmVEwDJ
slGXAL3rF/xz+MMceb4Ml5reDFU45cNDKEvlvXPGUZLiiOd/zUkg67OyaNdVuUQIf/rM29jhq/p1
D1oKLHfbjcp+EhrBD4wCB+ablVGhJeZ89fhJ90tVcSStsrEe7WnAiy1+pdUQc2ctVq7U8QUO9YjC
aSsWfWyh77rgPgzu2fGeuam/uHUiZi6prfxAHVE1r/DqC6cM/DFqBndmlahdU5E32/DrBMTRqU3U
MjXpkr0ONQQ4MIMIot/PaCoo+/MINIodB5whhUrWGRgLRnZaqviUBXvQfZDPYrQ5S+aUaxIjSnAT
6pQY2qzeY16yexEBSESDrPtqPdEOB+3b2ajLCGpB6JVz7WqGNDckI5fzf3p7o65aG6DGy+erGqoI
L9FpYOFQSHc22UiQ/B622xfr2+jjM9M/eiiTscbwXwYoLtzCuHpnf+oUpPV0X4vY1dI2w/WbJQ/n
16Wo8i2Gvn8X85bpSinv82T6rkExu7J0a9okHsAMNq8u+VihANnUD2r5F+VA8mTQQEE0yxw07TTX
mK69xXCa1RhqVF5tNmz3Cc1G7kAElDoE2pXND+XIojNRSKuMmZ5tycxYFhwmtabzCfjer3eDdQI/
EwwKcjaQkORnMa69+NqiOlj91X7yJVtoz7+cWfW9ZBXzPpZbTSo5/UMJO7O2xQBZHFszMcHH/YYj
c/oNLpjd/brAO91ORcPfm3izLEZnVPzAqp0oxlBr8KreWcVnU2k5stGzUmHZAO8ZAoK3ncsnaehD
BzFKrnZx4gj87f93+4faPfOb+qs8dsnCP5V7/wOexn4Ki5DbpSbC49OJWFRih6ALIIoWAxbLDzRD
67kmN3pmJ35qhXuO8DrL/ERrA2e1YAFfIq37PgMZhSMfK9EtaddzcnAHQ3inZfAMuJIqhpC0m5DQ
EKzvv3vm24XE+Eaq8+zvaTuRu3FCy3jDNt7HDOTViSxTsFiAMWrotAGN7fZtEfLAaso6yfcM5kr8
e9HZHcSRcZHvuJoHUfv8s3IP9vq6AZh0fTb4kb4OwpcwB0Auz2Uh7hfHWx0aS8voWyaU9DGX8bba
PFinzT9XAWOf6IWxBRFwZyP39MA/LMRgxU41O20U72IEBOXzkp5zgFj9dO5nP6eZMAaXI0lOUYT4
cXjqJFyBMHsgtHzWHozdOK03+raQSd8vkuFpQ5h6L0zBr4FSFW+sjUngitjrDZKtn8EUYDfUpt34
U1NzHeohWd1w2N5jj/1PLh2IHaYECtetYzgHSwYimuLN0vvgKg2rFAOpv2l5Iqc6WIMlGZSk7/SD
ZuDtyUTGhmqar+3RkJgSMfeq8BOX8doKnC5KIK16pCCbrSBYcweHqevAzZdspJHkQR3rX3HcQnr0
fZwbeNz2H8JTmY7clm4ABfuXil1fOmRRbsLamMT0ACA3Ws/hShdcPFsK1Ewlji/HHfZ6HAW1d6Xx
QT4H+AMdK5dE+put8hd+nhkdq0P21EWySkBYejCs3Ysqm6FNPrMtJ4r/TxVKQXNZBB2TAPJsHxQ+
h8V7hRJzqm2YIrGjaYAwRgo7aFFw1zQWN+RqR5prUOkn8snJRJP1CB0sXo9jm68/xYEnXjdtN2I/
mPF1auB78dY7BwBqbQOTkE1H/5fNjId8DDaJf44amuFRi689cLRkisdzo74kQDLF3mZFVjhDoeYS
NLJtiaqe7hAgjCOWYZRtUobN01IrtsokNd9TASlH/rETAPSLqmEcypyGyPOoEwoEjUczmwnQzhbn
Z2GXTzHFU6c777z5PyjJ5yyKUlCSt0zxnRCWyIY3YW1kvKq+Pd3C0TJ2Nib/SYVKEL5yLB2cY8Zr
4oEWCqoZw90ynv7Rp+JxHffdPZXz8a/iPk3CkNWfOdVDpsb7sEc15a+fhbvc5yzkVzOP5QHuVi1E
wGeOA8iwTQ/x7XLDIhh79LqpuDK0lTjWZ5xrrqk5oj0vkxvi1lhXf8MBoeyF7V3F1JhuSWJXmPKA
A1/RLLWhbJhTu3QncRPmP72Kl4MDGc8qKlxyiNlN/0UrU+Z1k57xzVgoQgibFYv+7q9yYS988mFs
Uy4WvoHD/iW78ANR1Atkz9UHCdP7RodppnSO8caKNxjEmlIJhHXHpVF2g4f1TrC9hGXH45l2Nr+J
bC4+F7aWbnXDbmCHxSg4kulkm+X02P2xV4zZw3LzIGREt1qde1rHB+n/RymPfuNK6ywfZbSIJjRB
akG5GaAYHKP8H0hGBB1C4nH/tvVk31S6fmsel+JR2pe7WXvNMWU9DnZWgD6Jwuuakq4PQ7lnBaaz
kImslkpM5i603Ohx1a4IxvVXBY8kfYDGpJ/8UIpvVZoCKMrSNisJEK42kAIAFcJCAYys3Wkd9LMx
VRef2jAMbGeVPbbPSWG1jbPVyHXK4iTc6JpuM+ToOQslM34TIhe8+U1Y2b1bu7K7NFnEv4t64jST
JxICZT4gd+52V2v93YITll4GbevLbHOz1zN+EwbgzRrTOum+LDcBpaMxn6OBGnwdKrf8b75gHgEt
2Kioo45BcsI9WdEj2l7UepIHA+3ngL9A9wcC1iod4VCPtLkrd1N4p6suHA54r48wEL+jfpuE5W2t
e0PPNZ4lBIMFiDbeLk4fG4wofow3jJW6BRYdBhkIugoglu39EWPARDy0ympQUqo4FoY9Ic8uIyK+
KNRfPHXswm5N5OCJiVVDwxcuroVkHq8xWz4wOwRy3AU95pCiOODgY4/OB0f0P5NtQ69/hISzCh/J
QvRDNN3dGob3Aex0jclTPrpJX0UnlS8Z4CHCuzzZ7EgH+5+QOtoJfYVhe/m7HcePynVHGInBjxGg
SxefXnrfIHbatu3fpEmLNHScxG/K6Vs0bduR1ls5kiGH0Hf3O9RPdhUW/hrvFiQ2Dq8tFWn8gKTz
baSoGEzPDTN4FcQJ842gyeWf/WhcVFkVujJ4EK3QEZpg3TuvFh/vn3mJCBZLiV1CQo2/D04rdRGd
IzOoQR22p7YnDgvYAEHDfar00vOyK9IqedbGwTibsraTsHjgAGt0QNJ1kmYbPQ3yz4vxUOzM8PFF
YasZthXbOMl8BDsDobVxAeuTCSz4BSuM3z20/kK+6Fb+EvVNGWFZJrDsx6KSc9yD/+ZqW049rx/Y
S4ozUbtJ4JubUkzgKUpebJvlRkTFQoWQ8MWs6/x+wvk4wipprJ8v4SczaZUioi30nzqFg0DIMJHa
TbeOIuVqmaxWgSbL6f00ybCmCyfAPMt3gOTW//6QMgGYgAMzYxwz/MfJHQfCU9E2JgqAvAWSy0eC
xthaxiKMlst0D9AvY55qU7xhLfMIUcJmIM0xpoEnNzJgQdMPF5SyqrWJUS2dz9iXHkWpTTwauO8X
zxGy962dxNSUHNSMa8bMj/WpwcKVFfkvNxVD37zPauC38jwDukVFhoNnD/XpeTlUJnrPtEdlZIru
kU4W7UySM/37TzEU1TVn0kx3wdAAOSbzeeZqsN6sH8UuQeShHJfQU57TT6yh2tR+sD7xfQXz25vP
Kgxr/EHIDaYP/c5v1dQeW14+aQY4rOHE0KuEVxq6lQ+MaZLg8yAlDPc8DQK8xFH6Q52yXVIOMKEm
2MEw9X+CINX0PzTvAOs9mrQqyT9pzOxwRCoD7moHhGkfX/D1IvoPjjSJRe46R1ej1TCmOUcM6EFP
xe5R/uv61X7fze5z1OoIfovo2LbXoT65/kjLtRMBu7TCaJIT7ZZoZu6qg/UK7V0ew40Bs6ghJPnc
UCai+Jm5NttUmJeSAqQqkJRzL/kBvMgRSO7x/hjC636k75cV/ZATHX9sJB3aieHFDlsjRL1J9OdV
YNCE5OlObhTTHJGGbk3bM5ZYrrE/xF4JIIMzRjexbhJdURNRN52ZU+Hqc0HDhshbidpJvIDXGi0/
klwrsrs+Zty9rbil6bS+PPpFG8lgvBB49NTM7tjBQzsGOS2gGktqK9s93DXyqi/wvmjTVeI8HME9
YG86bve3o163uwgs5iRzDK92xWkIJmLPBgvNAK3pEfCUXb5hceQf/U1KDyQktltaFTJZBdKr7PGp
l9UWTDFWZZDFF3bVvKY4dBc1epGwg7DH+MzSIDVv5HGTzLxqJVfH+g8SJ8Uo11pzyEc6NTJva2s9
ej1rVoLUqkkxDZdmOu75mwLtrFuQa6vpnsNxZD8Q+vd7aDuh80MmGdrXdLowiZw4Ee9Oa4iM2o3l
HmApcvOx/ZVUDOyqdzCSl/EFzOzDSHOzkRyPiy2cIFA6e4piOjDNi2CZu4RyCw6oafj05PN3AiuC
Rx9lM2SgXCkEHXAXVHgGSsO3YDASiCziakOP28GdoBbJSSHYWFU9AP6ICtuKGyC7QJebgdiN0evu
u9HFDJuM9JhbQ/1QKnWzDIhtOMMKyOf5mC/tslnULA8s6scThZOds8YhmLBKviR0T04ZluWKIRHI
2Dyg/kLj3FN8Ooo8yDqNHotalrYgMOL3nzw5xvdYVsIGj6ShPwn9/XeoSkqeku8WPyQ3tQIrGcfS
hnmf6Lac09ZBBA/bvy1gNoITErpoMzmkEABHf9hiNojGiPyx46snzYH6ZwnbadZmc2L/BCiVoojH
nUQYBxgY4t8HmnXUlfEokH2elRSnMIKRdAcTvSetcbo4FF16VaamBUZMsJN30EFL6Qtem/Abje0h
j5jHh3/aY4DjI7fbhrsUKlQgjUFy1dS2DiKgXyRA/SCs76ldS/8dG6e4kXTEp94c5Ox7jxg53Qyj
8GLBx7V7QFosKq5T053y6mbICZzCQNcG+6+6wwdotVZ+Msw9u99IR+zllhEpnCt5uceMmBgNHI61
MfMojbnyPQFfvlRigonvuiyJ7xIhw+qFeKptgCVaqrsQXJUgngo/YYiUEm50HLxfvvmGKizfX1Cu
H7GwkN9yTH1/+hkZB6P/ea46s4K1H4qTv2djspCwb1k7klcPiSf2diEsZ6Oi//SXGEgGsCoTv4+d
JyrhfJUnli5fKIEFG/7p75tv0blaknCwGEgsopGG7/Q2PDG/7HJSuR/LOpdyzAVraQNJwds6ETAr
emaKThoySGoYaiV3DxOymE7cMVOEImuDKFnUh6rSDI/53kLhpSj6MOL8ou56soyzSLGeMKS3BBl3
B6AzLFYDbu+is/LuaMburS3oJPkym1GwQ/FBzXWmjvrUt5y9d6gb38MByYgWjvTwVNHyKT41gUKy
GTXWhc+dHoAegiBvQjbdX7REpn4zhxzK8DoB9YachKHn5rzIleomoTtpwzo6cDaH1rRBf/TcyiGx
QFZRNY18RaS6zj7tettDQUY8IeeYn4MvihZ7Zlex4762p5+DD6MRmyB9mJhiqWoxxmU7k4Swxfd1
ZngXUynBhHRtecJZWvNm1vrZujH15wRo3Fy+6R1mSZwD6HuQ/8v+FRlzD6AHE+ESVBFtDz+/NZ5a
l3UqHZv5AlNWR9TajPvIm0vY7AFF1RTzDQsNxVB63hJqTK8JZV+eNRFDMxm/P4E8bu40ccQdIv1E
5OK1WFJJKgAYmWJx9GVvTlMGl5fPVAM8MXPGbjcznjY5GoZYJ+GFPAn54D8l8Uw7Et0gDJ/p1YFm
LoMwO7ABMcymSDYIj/Bxp5ZxijZc+LDkCwRkR3eTVFcisdQmZoM4gz56dcF462Nz+4Zpgk1KQX6+
fbd7CUIeY9o1Jus8TJ+xAOfJgVFUs3AYfNJC0OZtIk1gOE8QWDgbWASOrlZoDp7i0j1EbluZgLjo
SPK+fHWpK36/TJ5kD+F1mRIYfHswPFkzvHCpFznMuRVWY0rg8u1K7vJEKigHQQUxzsRqO/BWTsuB
igsRX+eL3QIcD/YZppc9ojVXr5nWvBsey8DScpsBkYv8DGY6/3L2I0/OpT65Inx5jLjugWsKCl4b
+r2pltnaoosUuLDqPJ7QtMWDKA+qNBWqR1PmS3WJv0P+EFOzDpErUyFL15onMJx49ccumoOlHapA
6J2tL4zLlR7Lc3Xmy5jNnctrbsvYCAEoQMtYp+/eJsmxGiRHQiAAaOesqSKvq84dPV5mtPslzt9n
ElwGHKrr6blveIoflNx048SGGa/YbNXulALnHKtdixPSvEk8pkw1sZ4hpN5NQSMge21V7+lyCf32
4SWzoxSVh1V4xmASKdkKtm+SiAixa9WBl2biIqI4XDP8N9sYMXjJzAHyq2xc4XmTXZg0/7Ix+f4R
s+SnU6bOOzVK1UIcId3yHHJ8kST987EYxWcV0t4ZqMg7HVYF6zvASSddyGPo11vLq+9qSOpuKAK6
7VD8DTJL7SbQseq47ViqgSZ0lb0iRzxYTKIoqi28+m0UVF0zgiocdA5he5DSMhLPPJ/5BL3/6ggM
DYfDX8FoUmgwmiWyXmN7kktbM8hs7I9ts/hUVKy6FWSZUkPZ0AEGgnzU2UbJMHtgXRLjgusCprJP
c5a5MSutfDYLbVTkCYazn2gE2pbZPXe7octbq+S2yR2wE3ZEic2A+1Y2R0gYwgZJCNGnUO8tc39o
m0EbD2vSuQQCcRDZOZ1g8cCqgjE7MLwRh/l1MXru0rMhseNrjIDSaTKJcgNrnCUaACmLPF+MEskd
txhFR5iVT60AB3dhlPR/4aeGSom2JyfPI5x57lNgCr6zmJyFaw09a5MSVqBnuo7uV1fvV8Dfd0s/
dVnXI0tFtPicmA5OtL7aBMqBq2Q70PUEkUjCDKERx7hnZ/GcijRZuEPb1UmOtXYjt80kW8SOZFNP
E3qJj0wjYhHhOKJaGnclpNuuDBYkIkfPCarlMU510TEkooKbcyTqyUQUSfZx4d/7gH2kbpYrc3K+
mxGiWkBDsFzLLP3iifozrY/EuPxGxtVoR0C07mqxOeKIcobQ3C9dNc5pzJFh2FXWkDI/Tc6mWd3F
kGtFX9oauKUoruvBTGiaFltPKKCOVyj/1dQwyMlNw6yua5FiVfWVI/MwAOYWI0ZD5tRmPVg8WO7H
0/V8QTvmK/d9N64xjmanITzvt2u0JRhw9ITyTw5as3QFgdhf91GFy+z7eS5uI5RkSGe3ZOdAfNb+
ww8ankZQ/i82rwcQpob4DzDUPWa2jP7SPDKl16kjlwfCfEzBrkc2wflp5pIavxrBiPRJNMJ8dRkR
bez29gmDUAU17Jr/bUyenn8yl3YGSLns+AnpR27Ghk/Jsro8o/jofqwdvJQG3LwG0KUz7Qfpb6tV
IW5pXRSTMhQ/urAQm46ajke4yJ/AXpVxafUfv10osnk/LDStE3aB/nD95cBzAB44pzANx5dvHZdj
NDWk+aBKdDg+TjYao1ziZD54pWH7MJez2SJZ/WtvTq98WfApM/gqA1eldqZjQ2Amr0faccqQvo7/
k5KwLdZc2EylzeeyG/IEmC5ipvq77e7NB7cZOdaH1B7hBSVXi87D+w5h+aktqxRY77vphRis6tkA
iU2HpTAn3IIk6q5Ivah0u1gddGJATopTm1KOOMzXQMskW+GV7fN9p5WOZScc604A2remwX0GRs/I
8EUJAjYzyatvaEYeQYTVAgfJuQ4CA6Uspl9N0pGkFaGpFi63/o/YEetlJjdpo9omsW2xtNIFRyM1
hQQHdkCOyxp/3JiqFcGHgHIceTT8uzVLuOjSXBgZSNWhD3qTUryaKoTxUep43HvRq77It4T/ghcA
JmxsLgQt6Fi3L6hPfAB1rs/UzXxu+OZOA81euugg3UCr6XzlcB7DR5CcFcOcD4i+1b8eFP07kKEn
G11spmJHF8vmCxecErDwl77fEHQRHdAbUAycqbH9Yjo4A6ybNBdbLrvv00MqBwbs7hGVoTM4RHqK
yjQNqE+oDsBvaHvg4EaUafuf2cyNxXV1IgGqMp0bz6CimqijgZ8Gne8cCK8/tWErAvu0aNKn89Ae
3/79nZT4UsjvZlLd2sipwPq7Z1srXt/lUaSTZQrTKMHvzceg/AfLACKIXhP/c8Li+QFAYLL472k2
CXyS2oEuI5XN6uHD9CIQMJf3/nbzjEnSk2DZ49cJJhrAA/RSsMynwJtBmELNPeEZnMqeARUmSw5o
BWrUPgbZBE1avEAd0pD+8WtqJFEHG2+WpeNggTNOu1uUczrNrcVZOVbRPbJfrZQWtIV4niMRGFwM
dZyu+CUuVTnq9uvomPCCP/fyLGYXBryghYiCXyAjOJ6P7GTxsQldtVjRk1CZwpqGLTCyKLdPohRa
+eCDK/o2OaJ4pyR1PIJLJKm93SQjBOrPf55xTZR2dSRhXaMMdYqGSTNo0c2B7gji1VQK4npvY234
N08MVwPkAw9iuD/5v0cjX5PkdHedTacb/QQYtrmJ0PsQcwbXdc4u7RS13TGV+asXV/h0dL0jJbO5
tNfWWp6G5wVAM7xe4aDDj5GH/QM8hWzTWd4oheG5aABAE1DXBu/RFwC3AKSekWfIdsLynQyVem+8
Uv66hQTqwcN2OQfD1971nl3JZsB9JNjV96UU93zqI9o8yAYLv1atMHGavnl7Ql3GJnoPY01f7aM5
gY9lY5x96ntwZlq0qeP1upIbyhEA/0Rryx85mulyCGGeWDI5xlrE6LWoW5EbsMPLQK+uzS1VOThg
Q8gefdlIlEiiSNTc0AqrluPi5rTqLGMoJwevwBTlsNNHeFIRTMn0egN/k3Qbf8B/ngStAe7opN5U
LV3I9wQ11FHv6xeoSRCfMVUHvo8QABaS0kYu9Kf/vv4LnMVWQyRbKBbsC2XndEUY5AIKbAsXm+Ng
QCYOVGokqb1X8319FIxFvFY2noxWjiQozadGxKRYKLm1yJlWprDhpQ7DL78Jl2L199jOUXUl7Yny
aphBKS9njrh/T2fV1dfErw2Otea50lPTbVbxEq48asVWB+0MywIOA5GjgVgK7WJXQTbyO8g518Fx
CXKqdMUH+kK3M6bv1GkEZXlOkPSdcnpPRLcXYCwZGoODEZdbNpebqSLZtSpeGIEkPl8wGD5Ckf8L
Cp5mVCd44g0yQ1u9qb0c/JLVUKjSASU/41NuWFYX2bBBeDkGBfuZxPaw0THrc0q22EcPSoeeRA2P
Y+B81FNFs/IdZ3O2xEz2iPTzCQDe0LWaod/N3O4qh+KUoeQwlXcYeG7uQqojtiV0H9JePAJQ3sDi
Wz5dEm/TDsSbz+i6D6/63u8GiNUqDHMQpwI61EY8zqF3SQg7uMVdrFQJUYJYnu9Wx5ErEQpLYKma
Pyouk5GAEJGHi2/2h6ZQIrbEEMkj8CnsZet4xV1ZXVUdzCcM0A6GloNKq/QwquGQwhbSM74X6zIF
Z8CkqiEP2sVHx1cSGwR2D0z2GSXOygAdsf9YQCoB32KigW8mJLfUuFEGTzSkbaX2s9PShHe3IstW
xfhVEj8UQuVgOYl5GfGRut92QUTHhzVKGInMINpqzBu0IRoKgrzzxD7QSxUEG+V0E85S5H+4UbPJ
qiNoZX5CgWmvDwIb9Jie60rcdEBfpVML8e9SiYEngOhcHC98t4AH1wS+RkfWX9dGAQM/5ggGsWw4
NnFehwD3m2hFlAFWPUwTHCkv3ezQvu9YRf70Bl2//cgEspcxhDbePbLqzo+OKjiLvJJe6pGSR0+D
6QPOFVYn/pSfvq5MuioHMI84FQEH3cKND7hCzUYrQW5lmb7VBwTL/ZUdOX3Ae/pyZEp9pFE33n9/
EiLdB3JqSIkv8Et2k4pa0dAjc7uwBah6dUBh+Jto9aJA0/l6nNcmvOHbghSMnNAQpJEYNP4VCMqj
Yh/ITj/VxqYZ+3KMBiQKc8+VJLg1og2G80ofhTxNb5WFIj9m9+73LiTmBGyOyG//IbtwXvwGgTXL
Sv82+pHWbBfOsxAbwGtrUkrCmh4vfSRdcJLa7xTDBF51aVo2g95qGlOMEtFBKJ325Fu/dox6UJeB
zvvr62Do1sw9o0JXIQ8riqXSyN2DeSS5h+1Ib/a35kgvBlNOMV/TssUCaU7BPzfhLhAbkMQAm9eu
WvKlgZp6PAw/YPrEl3toCrOqYTaD+Nh3CLYvLvu+g32qeGnUNHvdG2rGO+FEllAdEGtQBUW2VHQ2
CuPzb1aX9mm9ZRRfULkgIumUNLiO9hZi0QX9SnDMQYHT5rrNYHTiwyezA4HhcQPYA7nr7OOGcb7V
yENbe7+urCndHlhoXPlhGWow+bv48pck3K5R8kcc4VLKXaBJz3R1ltOWB2kJc116perUP2GcwGG8
JCNAx2YqJlgu11NNZVK0eRd7IRlMGphDniLCfidYuOBxSC/CpXBzdQPK4JoSfueN/E16bY1zjDQ1
RyQ3S9rdb1uOYVni2jNKxmXf93d+vgwzMTl/i2IVoRYZpW+VMF8mwOYjt7FzGib4pk3z3dG+eF90
2xFevSZ8zLtCGlJrFDnfZl+7oCvhFogBBKq10SuRUSQKSIr2EwHYmd4ZYfjXTq4Myav6luh28EI/
NTZkLJxyMpjnapbzjaYqQv9iOwSj23u9Mr0yNnpEeLlMlpadID7Gud/fMqOaK0ZflW5ebTGZ7nQj
Vf/gteUK2kOU+/UDWI9w4r/7mh/db8FvbFMlCQMqznYUyTMniOeFqFttLG7CR5F+4Uz5KUSkd9ZI
Wba4aD5PSCmMc/opz/wNPXPGD4svzQK8PjihIrY7b5KCCKTBd8b23gxKg7TH7BUtZ485GBXtzdpu
XGQZNCFbldAW/Ie2dbcydoECp+hmzWemIZW3vp3dkgg53GErijU+lbP7ApAAj/ouNww0cg0HBMv1
i6I35WYOPESPlpxpvJz5/wa02GOY6AClVXFp/p3rvTAdpkm1CqDkSJb68BGlIpjoOAkwF+6XChzB
J3542fcEiGZyEohFTdcBGpyuBeBuHH9pPhokFxL1Vx72o3zyHeCHZMnG2s2ANt/Z3lKR1Bplrl8L
6HLO0cmJhI1SQAMr2i+nTx/d+QHWLVc5zbqzRVy/Gjoy8J5WaysJ3P1FBtAStJ4R82Ulyam348I/
+3PWuAsY2vquyB6fblC3i7IgzI4ilZj1o9ptK0V3yjC/pBlo/2+V16Jl/gq1AezLYm2wGQMBLmD6
vCVh3zyQIrImmalxtR5fa1M8k/Sc7x7jg6D81V99gGH8Yj59jNPTN5+YIHOb1SuzwSYt6vhOVNT/
y6gJLEr5DZk3mxhG9w1LNw860WWeHUKCAcyYq6NvxGj5pxo7xd1LewOSSQm+3Byu1dZSTBiycMrP
va/mLu2s5Z9Bh8BWBuB08fRzIL6+LHeT+O0tZ9ddYgKPHGFDR0OOsqJkVcNlt0WcmLwMjvEbsigZ
vN9EAXRn8FW0mKUzP2te+OMRUchMi5QZ8Y+V95UYAup4dzAu89FZTPWiwArokK5HA026ReSrXjLc
c1hMeGVdWTkwtXszsYuVzaeTczKqLLYI4gRmxlshiI3+jPl2vKWr0/tufwjjdwQguFe09pm9yUSo
8UrgYqBlb0speD9i0DswKOYIU1pxsBN3yscq/BDBTOKFxlM6oIJv3MlnyV/x/rXiSGwr47YaRgJl
WG5aOasDlmPXkvxiSso9SZlWI8NzYbXGCwZBhhZ8nKeEmIxbZPOglv903Pp2l7XMBDjYhY+Fr6Ye
cXqXxOl7NUWl5U8h0OKTTRWBvXnX2/e0SONhmfosp+l7F5tpOuv/6xJoUhSxXz1eHr7eKMYyRmAi
mP24ITSRoRAfYy9kiEBKKyYJNiUMzCAEXmkBqnstEMlNG9XrylFqMWlZc74cbjPFuJWsrNKOm3e0
9ashyZHfDlga2B8bUa8tT0BM9n1otZVs+6/jyJ2Ob4z9/FBzBkHqe6wXbH73YLLiazE1puB+3M4+
kOmx7WPaFdMNMXelJZFQnvtG0g8WtZ3KerLhRGatPHlgMcntIXzqDyuYbnfSI3m+v3nmHS7hZ1B/
Z9o8Lx9QzoNuW5mVeyocYtrKVHaLawDtT9Ng10IAKffa+NjktIpjbtENEtJR4rNUVqe7Hp4ogJ/A
2+u3ahrJBTSzvASlDhuC9jwUnhX0Pa8r/0wXUUqcfoerFTTUwpYOS8CYfD3OGdW2Knk4otrtvALE
mJ2/sS5j09WTU6DG5KJz3CqYx3DWnMmDTSEjT6P14Sdzbp5mU7Qt0Pq6e9NYe8UOsYBQWuZbaQDv
nRrxZDmpyEWRMlVgjLPj2Tu8egNZyhHYwQuEJUVlDP9/ZdPgg/MbvKsLffk9nxu4z510RLMcWi9S
DKeh0uSZu0nQilJjurh4HJYFZcg6KeTtGXZ3VSdCpOEq/+SdnnELGvcGq/lfBhKo/xCT8NsmFANg
a3kbYeBU82rdaZEa33lMT8sXjZbDWHWSBrqJcNrCUaQH0bVmprvuC6xz91xD/cubEsgDWZxm5KcB
swpzNFyU3Q/Yt7D8n7TiN75fzyf9V8pRwa+vqC+pbimpYMlhyIEOH1EtDVtS8fiE69XFBUXXF7/+
4pdNBOudrr8L4T+nIuMPuBJPxyCMNwhEPwt/bJZgZEabqc1txUo7o9H1p/T/P//BE1imMWxKV5r1
cbz+Q9sQQ1fQjn7pCXXJPVR80T7OH0Fze4rvtU7b37dXETGYnv+Ua6+YO0i3d0qVAfcbMJDc6Fa4
rTTUlYWF3coJTirCCFsqXao8cf+zqMa12R+JYmKvBQXb6P3ajKXNUaqKaO/MPg5Wwv65fX9qYH9B
MpqBhkdt5VtSFvLjF45DtuuwOt8LgmeFV/9aa+y6mP/rIsbht/dhhcjmwzido4dfXMJfeqIk1Qwf
KNyaxw56hlgYOvgKUcXr9Mf8tj78OSqVnpJNdvB/9flv9yLoKUIbCnrGyJ6Yzoc9soTag+bGQx7I
z12WIvXrsBoosPDeBdKRaE5hz9Nw2vOVVd63Kyh5uHaZt9Os8C79L4QPC6udOu+taOGjLIMfUsTx
z7XPgXShzyhcdZS2NxOGsJY0fIxpbS1mr8rvJ3to3hqgUC/5BuoPDzuikCXiOTr2QUlLxaALnAco
MGHwtS7HLu9OSl2eSjRgsqPTA9bIks1Oj7ysl26bKdWHj9zhiHJmYPVxLd7s9AbsdEUg7fB9kTxT
dCe5iwRjPEr2ZpOEMbl05ZTkB492UiibBKs8iWk8TtP3BQahCd4bO2Tg61497W2r/SrpZeHSRVUk
pyxQFHxsibBflKtaa9V2+uQY5jX1cdylFaeB1ib+koy+DpZ4/m9msB4T4/7n/qSpIwMLKBks5gvh
EHBAK0/yJ89pdKbzzmewEH+3kBzW4Iwv24+C0s9iQemUtn5j8n4lrH0EL2nclk5CsQcWWmZmgQrL
P753KYZegFwo8huU+Hhop+hfWI0Lm39VyNV/BFcRa3BARCfzR7fGWZBuT3kLA0idzWZHzk+g5uAl
elJi9DkmueyMixNfpcTODBDAbrjJu7kU93u4AohMDrtsEkjcEvA8cIGDASGzdvM9adxszahXpEP+
DzY1JDDUMeLFd3SIYl0KeHgCNGNCavrBif3SjE1AcT3gmPahqwgosK+LrFImIE5/Rr5Sk+Br4WjB
gA1KNmF8WH32PP/WoKAyt2tJVPoyAZ2MgwMUKyJAHZvfTpXBopa94aaMUb83vTXsvWd1/k+9b44B
q3f8J3/OBjxuGSAf2e8vC7pvz1hKYdi/5frG8WA9alUdjIqtcPiyo2I0T+6MSf/rdvwp8SEYLR86
4Zc+nxLdntfwQxqRcDXc3u0MaKgdCay8sN7sRxc6rkx7iG+BhnvGuzn3a+wIzN1vAmGBarPmW/6Y
uwCjkJtfbqm3XlMeLAGmZy26axGb7h1JeS0x1skgDficHDDY8ShE+Kkr8Z1YPIQtS2bqwSqwHRUS
3/T/5gaxiSDU9tcYjGi9GYjdrSdMvLq5XLsu9qJW3J371tvXUwaWrSEpLdbB3WKXh3Jg5wKson9R
69WcPJfhYqOBlyUcLVtPBrxWviPDoOzZ3nfi5OFo2Z6j85VT3uxsHPc6jQMIxzR1DRHL3d7WEQNm
1Zw+l9fGMdiM62Uyq/PRDb9CFRrhmmBzqRCfcrhtKdHTApgSIOQHwzZR4uHkeWU14zWBVvnaQp/b
HsL93fBIr0rRG+iHpZyMLtY86eI0MjaIyVICrw12M0uD8UwfZDDqjJcNPuzhpI+0EP9lmFzfNWsy
bsonOSOlrfvVdhHJSLGSKWgQUX2yB78aLejqqCdWQEZiVI1dHo9r49aBLuABe/qUH6icvCJtzQiJ
gHcZHlwz5v+Bnh+JEGSd/M9FFuZ/ay01Vg8h2dLUAoFS0W1kX5FUh5iQQo9kLJ3NOF28AaU1Q8/g
si/7hRkRmdrSx4Cz5j51gjiPdqJ1ndw0aT5W9cf+AXk8x0MU03MlICTpF89KmJwOL6BPlLa8IxXy
Uk1UbaT5hsWaeocntrqWsaFP/f1dHdnj1gICkfMy7cc5VU7+iuwmtE00XQHw8GTJpDTNwF3XLHwE
O5HHkSz1+K6JcrP4tzpZGkPfdhoO5h/4I0fysFdQO1CDDTJF9w5hRxDOuW+7lqXCZ7sSGLykrdCR
xl1yEaJpibDBIq/J6CL+0K77lCfj41DxY3amxFnB3VycpFH4B7+zE8YfO2b7bRL6IQiGuQR78wJU
0HkbzXt5ftD7FQnHY1U4st6r3TX6BSJTEkchhdLBv4+pwk8+3HVz0OsZdXqLWanskAtYnsJIv4y5
rLAF063sfAFAo6ipbsrQvHAToxMdWqqtmnfXySlR8CI/HVMtp56jYKT8nRnZTZ3U9uBp0x6JutQw
ozuKzMpfnWgUsngIrk0VniAiMdhJjFSOgmN1jWl4/BbjmPlbFfF76L6cBIfejuqCF1fp/V/id/+R
mqRnFo63PZBgSxPatJQIJspfLzwiFB6on0KqR+9rwfOQb/QUrQJ2++/LRrLJo3feQ+eA6cySF1Bd
cJ9NiWpWpnu+53VD7Hh/+/RsRSIeehwtok6W25bZHZClJD/SFrKSpc+PEyCAFpEeq7mL/FmetiPq
8L/R+Aqe5j2je3hS6j+Aw6LNg9SSICj+IY4JRiwliSp4CfMez8YTIauOnXMnC2iFDXf/C3U5iXuB
vlUWWxa4p2ckLz/p+SIbTCs76kOFJqkp3oWlHQiWbksOC4WWJa+jpEug7qDxafoJlKCvAkxUePEj
fXHa80/hGl0be79UVtFH6UrvINYaBV9I4RjguHrTQuffx95wF1nW+AutH9AHTLixxnkKqjHEMl8M
+Z+euwWaNlktRheM/efpEplXzkm66LxpHRn7vn8e5CCII1cUEPM9hCVsQB35DWNiYoBqpXobtVta
7pnS3kh0JVCyXL/cloep0J68JW4X8juS88tF59CFWaQ7BY5yjx9mlj/gQhx4hvSM/CRkc215ul1y
5mzmugxuWRc7HywV1G4CvZ3eiwxIClC9u96f9OFENO1GJhQ6407ZIrYblW/yLkmVRTBU0btuURVz
zw2BroSHdyFZklpZz4yEYzp/FWdyLz2eTiy9XuFP2JShplh8W4TTky/ryjGVJ+qfw8HUhT0Z6JPf
i8nJLXrhf+uv1v1DyYpEuxphXsRLvyHpro4axpchEyMaVWbiU+vTVbot3/qNksdoBy9cHahcLLoz
/Wi4mtnE9K3QwjqUW3RGBuPJdtPfqPWo9AQSejHrSq9WQlzj+SgrBw3hBjGILTLlkWgr6ZHH5815
lofhpNJgeSHA+3xhglFAkFPeNNKLgHHH7QT/LWLvwCeJ46JJDBgT2DoHtWZdws2VyNFPknuxNx2k
m5Ajy20UPEJXq4ns86lzjZLm1ZUzf9Q1PHixgjGwfoj3tSZ+QpFHnfj603bQnvASy/zsNFrV79Ip
POmZRKbS0igPACLR59T/FShcrl7eLHxxfRj/ewggz2uEMXQjkuAv/qdZZGBGmUOi5RqxNApQlmLF
4BoL3hkLb245XbZBKonyBARIzltd6c7cqzSrP8dTPbi3+B96OXtzcvDQdHOh3rTCwfe2j0yogCX0
yzBtn6C8NufNmyFsQR/Pl9rORPy7K55JiTdkwY3TM+Q2QxuYseY5AXvPyzBdeBP22Mtxq6QtR+/V
F+2SKjACPZGXpM9kwHRjJuU/jpfEC5EfAyATfGmyONI/NnuW3cZSUSSQKwa3OtsXB9S1WhptkZ5K
6wl7imcTa7pncuLLMxEJ/A1mPjYppfsOCjq89dlBrdjK8N7cHgkTkWhT4zwnvDBdtbK2ZF89uzlq
PGFmQI72S/hyz4zbA1eVCQTsj+xSVz/XnE6h0sjgoHmkQiX3IU+5TCumlcuhe5yS5vXTFImVeyRx
PfR61es2fstfzf42lqjA3v7adtRNRzUasEYCfn+VlO58T5G11HHqHbGIlUKXJbqbst/NEudgTR2D
eDplUYlr/CCQm4xIxP9aosupZuF22giE9Gn6hOVx333uM0cK12rNBU31jueFtvBfkGz+dxkQVGkC
Hk5YQ5vm5BoCIILyiadiP8OQee0RNeYepuzOMvI19fkWB5lZcr4eNHPqgBcAnfkxAVl8IiQUeE1A
vcmMPxNIcQm/xQpsFGzDXX17okhYfd6x94SUyNrLP34gXBadPYiFgHnYoh6i53aeM5BCl4wb3sKQ
fDbWVlJQUdDjqXEAnaVAR0S3AkcUfYmGjZXQ5gMT6FqmOEx5Ot2fs2Z39rqwoa+DZ3V+nwy77qnj
MTaYaow8Y9vouRmW3gjVtG09e60kXbx7MzXg1VGxPYJVP0tqjDQz2BaVANEl+ZhleGr2H/ENkBQQ
4bas/hZt63UpnRglGOuiMj6/fpe0zF+k1scodSu3mggxEtuO8o23cY2l4f3sUJZGON+80V0oulE3
hGLZfjdU4Y8mh2leICAff8yMMd+u2fT+doTOfrHI07W6+sNaK2ys9oVWjL0AO26HLrMUqo8Pd8Mw
0EzXf2kkdQL0BTnEI+1a38W+uEVpq3HtgdUYkQAKv5rUggm4DBVmODmC2vVyHjOCqj8tFtuqDT0+
u7S8hbjBdbV21XkOUUGbg6H3T+T0JKGTIMMxDvC8po7LItyyPCOPCdLu+h5RMj3ip53aquUeyqrR
x4pA5xS2isUejWTzkmQnIby0zLKYzRiKNbAg+dmrRrTwG249qocxV9j1g0W/LTN2jJsBTQOg2tu3
iHKJgjDxzcHFt1RuPbt3dHxekSP2a0TqYQPCtj9NGnW2FAzPU75M6N3u4SBthXt+fNAMHRtwzhvc
3wm3Xl23rQG2Ms7OuChXK/wIGnLJf7+vmCSbf0w+nlWz5j5oLDH5LfC0Kj8y0h1+zgRBX1KKUm63
mMFS30+n/OOjm5JDRWXwJO3xvrkZRvhb+OlLXufsV75UKmE1l34eKf3TEe/c1qfC3IyY4gJq2x5f
0DEzonvBNULe4K2lE1zaphy4kb6s0AGXuKVSqjpjp9pmVwPJhnVQEkDfJII86OtNasaFg8lD62Y3
PfaT+EU0ZK5boh/OtUb2dt2Yt+YTK4cXf+4lYpcPOY8MWM92EiMTQ5704Llk3ecL1p9P6bhUEC8Z
0Of1XG0sU5jUMW/qeUesCCj5sY8UuV8/H4OU9N2G6vXvWlDgm4eIZLwYQh2HTzvyl0PFgPD/D1Qs
AK4BgEjGogqZdBiBlM2IxgwaJJRl3kap5m1WRMudQ0/4Pr+peBKj/nxXXQzdQceiM0Vliq9xjujg
ZNbouVYaj/JPzY2R/TKAY9PbxM2+WfW5zyZVHqCCDkiVb4NagLET12yJ3IRAK0mdQQyquNcOsBos
cVQWht3f92s5lTb1vXOezBw3NYdA3QlPE8Psn8yExhvJoC/eQ/PauhsDZGRn4bt5StXHVoqi0yQo
V49x0pHkBy+28Ks3lrjWp1PiYHq/EIdenngIDkWXIJaVJsJIUsp1889vRw9RSBuHXSUR+tWNlgN0
3MxeQsP9/CQU79Ax/RX9VGUa8eBhdXMpFqBdFIM7AkF/Acl4qJodW1+IZmlosk9O+cpT1yn/rbOP
40tr/3v8lFHoKDrsmNW9dEEQ8guQ5OGnGbEkKfxsMAkXI9WLmpiyaw7Qgt8Ygn69sUpMvQhEv/ID
tn/Tb+uwlKmJ9JjqKtsUGWf1zVQ0pIdTm/RBSivtef7DBbMXgp+tOBYplegv/AQ1InELo3i4mnpa
xmv5VXBNfIOgmCM0FR7nqU6ygwLlgmjdTmlB8+QmMcZ3Z7UWf5/LLrNhf20kDMjVgaj0YK8rSHqm
KHchv9O8MPG5cFDH4a6uGiKlnkVPyHkn4a+hvH3LB7IjqBafCVCS52lYlFbJJxzM9uZ7Y2j1kU+Q
fd7SNIPUQZGNoU1BXUYgs8yKCNcKyIenfUR8FvqhuEYG+NXgvblNAhqHPEa/HgFETK5zRM1IiIu3
/87w72I6y3eIgdaTj2mGoqf7s46R8SrN2W3Sm2qykThIlC8D7jVFr9pWrrmlISUTR75mChsTEwXp
rQcWdPRTEjJw3BrJ34aoyioQG5UanNHiRmMtDPnA291CaCxFOB2i7AQKv9HOVYZ+lYhLSchWhJwk
tTJvdGn61YFzit+HRz43+ytvlPI56cauG8jW3R7zsLjrUcMCnzBAAej+wZp/aT8DZB9S9JYeXtoU
4W0Ru7NGFgN/oNlR6t4RuH0Uqu7aGfCkal6VhRn2aPudgj6hU+lTGgs7jdmk4EYHYq/4WfZj7Vf8
35ueA048DKTob4K19koi4v0/THc5nT+SKTDIsckEjQRev/mtsie3a+KUt51gJjurfdGXcmsiUJMM
R7zCSvFJmCLBzOrLHwcmwBx+5lENbb0j1geipt007wlHgev7+FNZCDRbbXLAWtIoaVPbqo3YzhY1
Kw8aEOKFiR+hmctAyIwpTkHnv38gtrLbEu0MvyBeIjqiaPx1luytjjFYDf8LIdH+cPaOmJYMpIvz
1ArQPbNVQu2tKMEdCty8L6z67Y3vGTAmQPKyyT1it+YWPsoS2RKoUOeG62qIh8GjA8uHhr+7x3oy
Ty+KB2jSudv5+DR1SQss5XYmOOBcFv9+/ajWx80ekmkZS+5iaJpHZFa3sF8TNYZAgE+ItkXohKKa
oXqhTAsG+z5M/9VTahnLlzgyNiyNxH03q5536HTQOOtPG0mSDlkL5punQxoUOmOrEEpWCasIOf+S
BPdHwCtvjCqrJ/wdHvTR0gVznArOn2LMkNT/QaIUqAEl2BUe1LYpmeLyPI1z638O7AVGSuFY1OTu
EAphx+gJm77xRCkArZJPwhzEaTVyTgjcq2kta6ZKGTQwM5+PynGbWYUl50Iuzk920buTujXgHf2i
attoQEBH/G55E8QFYrm0rIZjH5sUi1438t5tIXU5c8tkBykkiYq96XqIVAtwYlSsul/IMYHmcwzP
n+09V/HZhLUoFUC+tzxEDVl23w6zlHUqCQ7zK0zWwG879Sxxx0GdwuC+jqjccHBf359LWH7XYmxK
7mPHCVWr1DkkOuC4xmSinUcN48e0vUEsaMRX5HydwjAUt8CmiRtBjnfi1QOLaggwoBdKhkPTz4kJ
OT4vLf6JMf3vKyCfLYq1Bh/u0RaW40sxtaaOpWjhqbeYgE86Qi8l7yOaRstlrz3azw38lJ04fwO3
rZiS/Phh3G4vaF6u5bmkI0F7ygod7tFXJZJc9KineMSGtsmJSJOa9HePeTRDMY/j6jXcr0HUI2Bx
GqEyRpKrbbnxcXezdLxIHozOhuBCz39G+7oH6MiglgorrelTgNmvLtn4vnYLgriDnzBdW0LRAfeB
Vb/fqTczFQ+C0yJpzTz1DgKmy0IF1wTt4WUOrbqUQ8ZTOZAVXIwXNmqv/mTZIPmKqbmUM+vM17w/
ieSB4TbCrJdTOYNzZr3apEXqYWJnp/VceY6BfRSsP9pWfnyD1doZvUJntlkJadidlfcedX6VbIoR
oqy7BDUoYJWOX/A9MUw447Qff7IQKW+b/89tfbeOszZ9vLPNnEh4pBbVWpIwBMc/VTAse9fqlyHN
Mh9d5dRsIRddMkxHapCMeR0TgdPOzBK2LZ1S7e717AD5wkSc5b4Xg9p/aKJmqqcBA8gfZJOqLmyC
AU2u/fKUX8lbiOymP9hzk3pzckBT6P7ap/GvBNbGwS/mdYaJUjgvFjnZhUYYfZBfl1Nyg/sPsXsi
j119TcoFdu9Gd4wK6FWVNOnTpbTUpAW2IePs5Dwene/EEUDDpAdpo+HsPJjBhjB+9J41eet3Nom7
Mxu9Z2hJfeKGxnasrwScgV3cXxlvrFDhVgAX43O4kOacSwFdruUODGWk4z91S3gnTUb8v7zwUTjv
JvLOLOrNyfYn/GU7kXUBE4udmzt40t4nGmx02N9doZuou7cSRSNwtSYvuu5o/NqOUFIS2eChkghj
ftmdyJSf9p0+dgH+ORmOqFkV75473a/o4UepuUxLshJCv2fhFbWv43CCpSTCXfxHKUeTsywPJYye
0YFr/Ls0kcu19GQccicMbrmk3i39M53ct6QBo2jyNIR18DzZgZx58iIO08qWcVLUwpM5tjHz5B+o
It9KJnf8txPl4nWIOR1RunDBtgUU7k/yUzav+7vv6WFOtWVS0hDJn/bA8jdDAD7GvMqWuo8BzBbz
dyBL4UZJJBLcem8S/B9GE3hBYmnQ5xzkC7rdmjrbwsg1bfEGNVFsFJJAlTXF69uil4oNOB9BWFiM
fBpgyDebLfLPaGQ5C+RPo4vbtF0w4wrspRUnZqXezAo5AZyeDyhJDSOQYzhJxu0ewZQxyuG4m70d
f5osFYV4NHmdrsLJqMguwuyjiiiX3BcGJ7a+bUiZOgS6//DVdJUZUhRCQuVjTX5jnf2at8ESKOwn
e5d4pbfOykAbDNWuSzeQPL0xmWzrZH85I9arjRuk0Bv5ddB6jwPaYw31RDjuJ614Aj+YgkM9zpkS
wKrr12+FQUXSMCLGWN7Hp24eQmPq01Eg9MdXP3LlM9SQmsoxW1AKM0z03dHjefBUfcIKC6z9nlxi
MJYo/LK5AvvIP+QQ+Afe40el3R9lnRfZqMErkWRWN8+KjZsUTpHRCRHLPZdla/LAZ4Jg+R6262E3
GEfL4aWtrCH39bfDVaObg73SPNWPvkt6d+BKJX0vwa4WofWkPvUeoRLBjRMIqf9Q8WOiD7SKZvhF
DQa+oPNneU4Ul0Cqythmfk7lyST0fP0Blp9RwT5tybJdl9FC5UqeX8GGVaw2aoq5UoFpCUcP8uTG
aqI+Lql2XHQlNB1Ov7X8GvuUWTvnHdk2/Kv6kgm1AHfWq0j753/JPptJQCzdwUzucYQiUFwUcTDh
Bai4JNzQLxk9vpm2EPA8joRYSTj+yCjguAexTPN4WM1TGLDgfAKLH6cV6unqiOOkG/3AYhhME18M
OLjK+Xu2KnLDcky0m0zXAyiOJP490ppR9nMYq+j7P0tf1haAI1IMXTaRQBtzMXsqkcvRw2sDkL6S
kCsX04nIuU2903mcN1cGLscKuWjQ6JovCN54qr7QlReOUMs60jkHyYIPLg46yMV7S+KPp8J7dSan
gLkZBkfKYJf/m9LEY0KotoOWHPe3N3ouUxx0p5+ZlfyvEBC2wysx4++hXfo/AEop3B/OQROG0m0n
CODVCbzOxSpXc6xCVr1xo1zbfDbtYJyFqNbp5A1xAMylqelN5HXCXfE9GOkS8JzAW5Jms7ATOtgc
WQvCZNJeAeQrtI7hHq784NDCPr5sE9VuWOEwFpf1PDumrlbHPPpBlOFNnULR7gF8ujX0YDIuPw59
1i+5ScQKMu4hsOFSNuk/ODBRGPTqTCbMafBwqRt6qHfRQyD9Zr6DdBR6BC+TzaM7FWvVRqKkg3kN
8itQ1yv9AlzWShZa80RGuZETAjX9MuBE0PXn5kUOkiDt5YwsoShnU3hfDJk3dNDm0zBdfKqg2jbl
Pz1Kroe8VXzddfHBdCGK/v9o8p6rEXI87yWZiCkzcSmt+Tx2o98LEjHlNUrWvbapxTQ74HUgccA6
Zis9BB7H/O9c+Oi4CuteZiDCV1XbN2M2EuMAb1GnFxN78UCjwMpmNz9NfxzAAxCc7SWitBi86R9D
OyNPY/hThsxFRjxIeuuNUogi3Rh1RyGgBjn61IHOfwhpvyYGqyUYhAgQStRtCdhSw86m+IraJ1Qg
vJIPLTqjE5cm0yNlgR/udL2KJgLSzD7tw8HfeKPeCebZ6s7yebsmLz4e9yQq6uGEa3YBdI6ju+dY
uEqfdD0bDr+vvHa+pjCuUrR0ZZVP2Z2jSwU57J6KBlV9grBYcycj7iLQMbpEtRMZH9Td7XNpXFt6
aPa4gpnjyfit+8nD+Z6QeTtIC6IgLKIsB1TjXRywtqOjigz2jNfmXjjNc3GHLyCbngyzJlKP17SW
P8DgUCjaURFgCo2NkpE3phOauifCPgLzd8/LIYP3mC3r0VsPuh5KBeqFXJpXy6PCpMtcX6PRcBbf
Vq82nVBxwPdbueYCnlAbKNgYXtUlwASMSRQgzw1pBEvTCxAi5PaYQ5Ezs5Zn0Bmrb9U/IOpZVc9o
70cosrO7c3gT1xLvWmn2GIvbRrt1twirnPmU0vKxymEByMfs5+KpOcSLrfLjn53wks6Fc9LHmIyf
Gy3UnIOmB/CFMH3BuQ5A8oLp0B1+MlR3wn7pnUpJ54UxALgo0g5QwgXE9KH7rEG6VvRtNLkZTB43
HaivV5T4qY78qtVCJwj1nsE3C27cuza6pFcrGuJiD6a5MEM9glHVQdng7ahKvf7goT2ofXQws0YV
wr48hVPWk1OpyU8dTEAA8KjGxvVxLGHyvHqncdCCmA6T+YPxtzfvQEcp/yN/+4BgNBJhdgYy7ppx
isj9DVmCrXkiPe4nwm4fAMoAbCLu04Cpx+OOBCWN+rHgkitisVsfgAQYN6dKRhqT7tBI2r9wdvOK
GK1XWLrMm8IQPgCyCLy2LFEpWFu8BbIAiKJLwRqAps/RxRsIUirgf/v/vq0PU+X9zxvBKA7wgMyB
QbfjdR4Ze8/BpLA2RcdCT0+6Wdpukh5ig2xrZtRfC3NgsXowMlxCHn94AGSBMl7Xwc0SGfB750xp
XafHcVNgg3rZ6l9Yu6vCL9l/4l7velmTZjYwI2bMR2kctpnOPuaI4UEjhSJzHBzCzmrhxi090/Jm
CdxOWkESRiriGEUIggHIkEjaSyEZAEfBkFydmNHEvcK0IT1RNKfLd3MTACSZauqG97PToQM0lY5s
Uq8Jx1plAoIv5EBG2L12u5Em2h/EXZ8VwYnqKtKbo/jsUyWwKqizhFXnIEjDErh21poBLfwxcO3y
zsJ6I8ClTIw7ZAVXTuNRjnj2fEyA479N1Qyoc6xCa0T0vPWaPJTRoWBRInMwwJf5EESMtkjPV56w
DpuwzeWGmPtBTyuaQEqxXuQ89JmunUTNiNUS7yforfYVzvq0nZtbAe7uCICWtz7HSRtwGK5xtAiN
T0Nvb4BeO8qiUFGwBhhrCLYO8RqVSWXtt4SqwiFDuRkcAY0sSDd0Zly659rpHACJphkOqRn/M4mG
ACyBIdG28F8hHUqV62svVouIPNdpDPWqVkss3fjpVUy17hsUsB6kQ0cRqkCd9ys5TXvc5pQcHDBw
07nLP5Wfm9BS8o73F4fnDeHFpaXr0QlRddeNjYzVXaQxURRilEjDAwD7EoY+7yRwZOwRBE0LJrej
6f1WzZ07yUHsVU/ZHJVlWLUpxQtciJMekkhzvVy+GbVQcaia80ylSx6zc7s14V3Ht2MgqXrIv0lz
V7RBjJ01ciLzorIaHT6dMc5PdWyfE8aYxc8kFzTL+R/o67VWKTJujnFKCs1YlXlNATpBbfNZ8dkQ
R+yNlgIO0GWkQxjRJUkp/nY1Y2pwDA/Nrpnz3AzLFBGf9CMIDIICniot3H5thpSanCYKlNXbHKjS
XB6mr/LUd3+y6V/1KaLgXK10hsW2qcULk+bcbQpueeC7gSYc9xGpn7TjN6GZ13MSu6f31TDuqFJD
R3JQAu5y8ReiiOFujPlylUovleMMWzSCPwBF67ayqEOv2jyCW8pTqvbmAJd2/bMfhCW5WB5QxCBk
zjAq2/053Bx3bc9pq+d/08wD5OheER78MkUb4FYt+g/mz7YEi0wpRCJkoqRw7s5e1VfGGXHK6cfd
6gJ1ZNq+6rSAbtk8cO4bwZbNoeo/zHEojJprRZMHf7g0xwRmWlFS2yApvA9Q1Nh2wHzBp+j8QWAT
CgjElto/vdLc0PIka0pccVV9dQMSRQ8U9DG4zf7f+YlAXTSEfRAPGQJi/0JHeEtBrowftA3WEdI4
PUo8iSe8q3/KQbRtPtdKSx+q999Ye0GyqwW/GbPjBJy/g8ZO10UrgjukeMoD6gAovh8ehKQPzl40
BUxiPLIZpHb4ucmQ0Cu0jBb0DjKxd0qwENq7yncJWNt7ovpqdjzbDgS39pjNNKcsFpU0nJFIO4O1
rP8VLFPXlOpXF73904oQ5DPMmNb6H5iLYEIF9C/cKYHCZhS+/tYyO3R4WdrTUi4UCHDO0rk3jEmZ
qkOTJLhOdC4D8HNkQfBUsvO7ajRhpdoQaJuPeT5AwvR+LQ4HgNurpE0jGdzIshIRNyFqHeDH/XDt
G1WmWTopTTG8eDIs0fSjchDZQjW2ChUumb2dWiS6WwNzQvMzGR9UAeBYSHimlrzuvhRc2rdytczt
eBFS/F/gTYhaetLsCYc4R7RmtLzepqvtgrBQleRrMbPQoiftTC7hmYeCZ5ait/59Pw3EqsEq4J95
1MAWCQRpVdq2EPYaZZbCvisMtgJ1MTE6tpZydXs6jxGPIsp2Mx6n7HqqIrLAHRYbO5AjGLRq07lj
KJLsy09QSwZTMb6fMz1uQYMXOZtExnu/oT0+mJGGEZNFotL1cMyTPFYl0jy97NHs5Q9PfHqck+4U
mH/Vx/XQUG2/mrNMGFzHOtso5xQd+uoMgSD41Q2188hMJTBw/vOzounFOQgGO8IMddIri1bncBRW
zEqpTt0jNwsPWHi1vcpMUD/KDE9S43NxGUfRLYlB8WhPDhm8+MwyKM3LPTzUFpFhclzLFIjm7cMc
d+kJl/vBa7XnNuf3duQma9xlswRP/mM+3pZuBPWCawca54yG3HUmHAJr1AlbcDV0vGis7zC7LamS
OPr+lB99Y+C8qGOIq8U5fOtiwk69M0UuWMl4p7Nkzo1eSzoef+SPp0NjWSNMDCJXdReO6U1wnerE
fqmjnoxgL8jp2N2Pz1wbngZ/bWpBIhI5pyn1ZCmyJItiQRAR816VxvE/7sdLpObErSBEgG3jj7t5
+ETbV2gfePVBQgUnfW5MwST1qppMPK4rS+okLJKQJ7WGZWgwZd2OgQg1KeRLVJ6Q+vcEK/mvaFZf
2cyPRsix7uIG+L9dBYTbYz431YAkSnVwJya8OQbIeyhHGzTKzQ/t7f0fpAd0XfTJQwQijtoFmlSE
RT49iwFtdScgDSI5q3eme9KVrZzTn6Jp3PuRcxvrkmcpJjgo1F4eqhLiScqmyWD4OWguzWdzXF5X
2layDpaJeCA60fa9W9KL3m1Er6v5+pthwTDs9dwAsmRUN4uSJ63TV72nCTsdNocLWLc739hMXHOM
xNCc44y0loRYEhRnEM+OG0g9UvfjBfLKtapVWUSyA7pwNaycqAdTV7RHzsWzaZlZMvbwGtSTps4s
HzbMzOK21K4Q+V6sQa+0fIHo3t3w+kDbnU5nrPJHSh+ob6z9IMLa6Wypgk7f3/9RG7uSDhtvGdHN
3K5+gX7vQtvkShFIu2zCpxsDvKA6V4or3UYpXEPv1s6RzUs8xhDwzlyKBI7WQuP+Y/sxVd9WFlva
w0GfkhCVdnGRrdzDn7cu0G9UbvhfJ+FmDKcqvxQIUWxYilWn4JLpf+3O9LoYrUwdsXxIqpzihiom
W7U3VDNccY5ozk/27ob439lK7kvcYLW+jUlwrKxT3JD4YNWtSjkSSayWaUa3cVURAkldLqtrt0ia
C5ytnCct8qZpQF+2coHtSSXmuXovs+2nptJr02nF33lcHY49ZHT/ViHZ2MjK8RmqCqxSg2se8+wQ
VXLHGReraJ2QQmSLse1QhiNNa0gyCMHfEHOMZ7M+lm1x1f1kW5RMShBjufdg0crT6Wr2MTq6OHuU
PxU6PxHExsJdcjT3DPMRk6WNmnT23knqCbR+s3QRfvsTAgK4VIsmAfm1FRWFxN5PlBdFRvYX886d
2wLIdmE/JQk+LuWwqiGTUEYv45ZMybafsx/pXx/SYE5/17I1xPShoc4hFchVbmhRPoMWBIJhvzE7
ArnRQ1uQ1Le5Ly/tUgAuIw5YllLp+nGRT2D0ZIn+pFslvp+aU5fpIwTOR2u7tG+z6Yq4AmpGe8Zh
h/moxaYvzs37OFEFEfx5u4E1amUWuvsmOMIRicgbxMnqoiY2PJso/wPUGzYnLkz1262J9NyHR7d4
a4e+9BDL/Rzeov5qdDtvmPGlOqkVNjtRBxxFxibEQOfHD0+uFUFr7dECFSDpd8w4JRno6L8w7vAz
SMen5SJAoM2tt48nLeZIzN8OwFG4Leetg5LuJL+0ez3s3lagoR0Nk56LK2aV8NSTyQYIOq1juWGv
QaaJzs5rY+DeKILl9Hr6IFpXM41flG4wIcvESXNIe7o94/N+GcBo/8+jOGDvSxvxVkboYXUevUMk
Ysyd0B10usSmySEmWKvIZ7TeTbrBHBKUcBptqCnF8oEu9Oo6e4zMUR8iU5qLgbksPW0le1ou+JUt
JTkILSCIYs0msOnLHWts6AzH9z1679Il0zIpaHvLS+wLg7oeAjGR6BdP5VPmrXe3w6DYiCkdZoAJ
xq4qHkNbR3LxnWU2LolOndqLEh6AbBZ/Bqqvfw7Brp/Icdse9WvIjL5iUiF0HL8UzttrU5jnD/j+
WjPqhERck1rCADd1YWP4fN8BmU6MtyJUG8AiDelM4mlML4ubhKp7YqmDqawBp6GLO6IhQYwOzXNH
KZRG0hdYzkxz/XHG4fGFx0f/lb/DHHeRZk7eXs5MPUo/AD5EuKReugBavIguDMsQL64g2WhteWPn
C7TLD9iuZNG3sO7CwA41OBRhuQqftm2rCydxft8AblMLWdztbo657mQ91oyaTYqpTQIinZs2V2nI
kouqnlB+3k+3OraoV9Sr4d+QEZ23i53uCvXNF7yXd2bf7/54i3kTUfx1OayXHIjnCRCH/yzisYK8
qA8hUw4dG1AW/cAbGljXKP3pClYI7SJ7kF5QeZ9gxgxkdhlJ3Ytm4/CJZ1BRaEHPHd6GMWsyJD+I
p2jIhoEofZEg3T21hCG/ddvKQqaaNcXICwkiXEJ5evb4mwD8TNFgXGkAbkhDzUzlDHF1kw+dTSr6
TlDbZCKzc9TpsJm/4sjo3fXWiwnCZgCIrcpRe85+9AxvwedtxAn/hZ2MMKYPn1BWtOJP6FYW7HCI
eJg9H5KUpruL1ke5xQhmlpUSVhMZBQIBWbYzGgjV+HkUEcCfUPntIHz0OUZ8K1iDW7b3eHoYnH4J
NlMAvS1g2IfDiWFBzRKgGj6bgFCqaZjOyxO2i8HaEaV3Lt/D8KIM+2NqK6DSbSorqhWcB/6DcaJV
w3+nWS7sl1ZgFiE1Xpje3ItAdySPkKQy0+03Gs2q9gUL7TTMHYP1aEoca1Ehghfq3qmZqgEt0KrE
Exo0sq3wak6XtJmhwCjzRrpXtqQxraFTBzaPVOSdDOFt68pyYZ8L3LgHRndZc49/K2DPKTtYKa6L
GXyNeUe0ydQuL79pEXQTZ62ISX7ZhY03W3ZamY5Hy8TNy87gBykIVTFsBxjeBXNw4C+yyoANykxO
fFamQAtiiHMcMKHcrubNhmryUr/M6VNX6DwLFOJTZmikF8xK+wK0/BO9DsiaFHWhypG0YMvJmy7s
J8pBEGT8ZB9ozY66iX9C4xKUTzMucMjhXiNncB6qFS99lH2gFEDupYDFUnCR1sAWqObPlG47yN1W
IC4dUZmzAXEmQHHCHYPFSGVhOuEFNPuudvC8KWHrzZi151cAMIw0nWhuyzUW9gPL5lg70g+F317e
zWXaM5NPknX0Sh8s5oSPTm2Yp3CF0p+ugcBKie2QuE3N+4tdKZAe09YAeuV10vcjQI1DA5IXZRxO
Wy1OMHzN2MLqgdiv2OiaClLqLYhQPUZJd3uN/sAy3wsyjHTFn+M9WGHEo4450GpC9UzhebCG7AIE
WBT9j8plkh4+ib8yG2d7MfYEY0VhA+lMVA8BI809pYSkAik8W9J8AH6jEpOiewoF0VZhSJCZ4aUQ
3R6iS0OVzP2IwbdI+i+MoTxluM1qgYE0Z0M7Rm4eo6ET+uV+WoxpGNPHofwR2GjkvKe6nLDbC9R/
Yp1ItehV2bTHqd2xz0rn4ougCMMGQPsU2g3kGe5simIU+D8qnsTIjoEl+Ssrr9eN5qTHOCrwVlmr
4Wbv2UovA28MmpXrpuoQiRlHY8T8YafF9FMMW9Z5uYQcgeBmfCL3ROb75/4kmUyrhj8d4bge4xzx
YCYTW+TW4ZgaBukzQ7AQnSzXd/6X24xkmYDPmXH9BubV5BBHHdSkb7zcK7WfSHnAKCTejaZ34FvO
qsBVPlmZPhUqR30/bTG7IIaV2rTI1u9+wxKswzZ6kd/xOA/L+c08uBhtPTIQxRaIXK8aFqnBWMe/
owFcioIWnB9KJ6kGjhH9Smlb+mMeiw1xFWHmJUCPwGZCUXpGehsziCORRpqDTuVMjuztfnOZZe2M
yZLAAGslEyh1eWlf+woExMG6yIu7NuVnHie2TqHei0U/eiyx0oboN4gfe+lZ+c8D085cfFWG5aQY
oPyepvgdXWSksxBe7KrKlkETbxX8jaeTZn/tpkN0QLcL7QgiDEKhrWWfReudrBpbGOUWSEcM8jin
YFVaviQmo4g/+blRIm/sJkQh66FUrTDERyKln2WpPtlIJ41EucAr/Q59eVujszZCR9p81zWHnBAV
qujGi7jPCza4hk++a6dHBtJoCLhjwqscuizsi8RHQWRMDNHpdeGC7O7C2d2VDkGyjO+xcbTWYDAr
zuA877q7Tx2XyOIie4w71EXiJ15dY77ovmF2oFXatrRkRDlsf0JudrDFCaMNIUQgtJsTODu+IQf2
j1/79K/k2R+Bs0l/sojtryGhlCY6NM0O09N1/3dJF207XL5HXwUJcV7a2d9OZndE/qhSwhaPQWuB
vvgO1QeCtzRG30q8PYc/P2JokHqPBKASM/iWVbru0YMVKP5dLGSfUSDnUhwoyKsQ2gN7MnlHM5wq
l/g8ZAuuKLGjqEQu1FD/L8scXBbsiaXI7F6BGqg+9sTYyfrRbv6udf26crXvUcQpAo5A+YGxUsSG
AG+i+tzm7hRjIJCon0MWTDTSxFcfDjRygxQoCe2R722zCZe+3HRy4Xygnv6il0s2/wGLp60tDjjp
/33t4fp4Zu/ya8Dw06MW0EiJ1wa0V6KNFLpLKwV7QbJQWaw9Wg6K+qqO3QeKAUD2v/K+68ds2To2
AzOT7xCGJjWwB0t5TtXIohX7YnwimcDERijtrESy2qDqlrOqNOWD6Gu4cza2cCEmTyD+rocsQ3GT
T08vNuQiDwZCFIDgyhnNnItMlrDqTp2ZPlCPap1E8uD8PNWu34WjFfGi826cZENXgfRLv1uRwUHm
rovJ1TXo1XpUSd+NF7CLAmJiMwk5hy99xd/Tb1GZIAjuQL2/02NXpJAJ3bO2QzejkvPnoUNoZGnb
54ivijZX0TQFMGQ0ZnulCcDAsTNl5VL1fH+8yvyDEmMD6ZpkgDkKkEtdJ0Ek5r2yBKPVELaWv0Sw
8cQ0JUcssT15u3t020vbKIMhp6TUILMsid/YaYVGrteYULuCCM/opGnT7O/R9urmqJWqPyZf9Z8R
o0H45mBtCtX/8cYSRnoJHHskO7Regy28FTLB8UXPZY+7wXtdsrGUJSgN5nS/Eqhn5ks6IAwGpbJy
TS0FlV4DORDvZL15lD/zoIMKvOYqMtwzFdxffvDn06G2me2kfiPBlsbxv6WxQ2rG/5pnjr8Y8PoQ
clDx54zW2gmODXixunHtPNTa1+uLSWsdnkpT2kA+2oVq4Bf3eC3VgKmW7c0x8zCcxJ0pnbDJ7JE6
TweZNQKrAo/iNR66pzEuPeofJ3Z9Fd2HsXbb6POxGFbByZa+RRoITPK3VWpoB0Zv3aCiH3y08v2+
6XZnAJqj+cI+Hn4tbjDsKjY+JTwNPySROgan9WL3+z2HbVIvxZI1ZKCbuFedJMKlL07YdKg8TiZm
jkJ/rDHTJs5FfrciwOn7r71Yms5IgPGjJHFUBKbQZaWo8Hbx7GuJrMrnG8AK/pKULJcnCGsVqyn1
qLDxqBuCUTY2ujqb0Ub+J1aowq/Mu8kW17hq3iZUppuk6lQB/cY6ORv+pGm/3eR5E6PUBqiO10j8
L5Z3jJU+NoEYQ48SBa9e42d1nxjO28m4jFOEAA86fK5JQNn8pKmittpGxhE9bsDq5XY4laP33OKG
scbk9UL6fN5hvdPAB9KQ5tk+UDk0EdzbjkYQEXATkKH2v1yL3GjpYvrYhdXewscqEHXOdAFljhmn
U4nRIek7382oxvDTVU3XE7uNBEQPH8w1+XC1q+XC68d2pRH5zPpsrv/ftlyE2R2l2ZbNxNpXJoMQ
IfhJEmDNP0z3DdmRjkD2kkqOoPo+iLKGEO7JOmiAsg2zXUaIXV9sHViQq5oWUZ9Yxbmvae11XniA
qhNXBMXg/8WX1UE8LgA7JmlxLdDPUneFRTYnVaPZVQUuCpwBiLcWUdVyDtU8IDz7h6r2xV9A049+
NBtGluI1LZICGVqbqupaWbgaMPszCbIpKWuejPo29JDBjOZuTZm/sJmDv1VUeGTiPI3bEs6OdtoI
XbzpCyIaRdUWe6/oKl6Q0uXfBB8bz0mW2LA1B1YrATXrT/a7/E8cggNLzv8BR3YRXA2ROgnUIaZy
IpQZ44bwGcpNt46weg9yC/ew7bDjE7HR9DIQIPhZ29VljnICdFwKnl+Lb3LwCR+paMNSp0A5GgQt
lUh7tyROhWc4y4TYWjd25F+xDzBXztqMhIHmRM8glCUKe+/pzjBI1vzzjPGO6nLeOmkAXJZovw9m
zrbo039kSqqp9QEWKXYGycmXa7QnZs0btC40ZbaZp1jF604V3bu87WN5WgmGwRlnAvCH6zyNeCzh
zziosS7LGuViSThmaa/NqofM9toSidapn7lUdHrREK/kJvdK5IFTN0y4hvvt7kLTxuYkyOAHNqX4
3ooC+Glc9auNYvs1aovgj7/hORXznMHi65hvK4KTMhiBGEVERDfOp1l0VNcojY5LL9ctDZTfIEu9
3K33rJmSGR3Ek9vZnGyrRx4Qtz1kc+T2u2ieztSjcN2IMhx3zDZXqZ0wMGbDJxALIVPUXThnPv9R
fAddKivdD7z21TMZpNJtfavDkmaFsBivGoMZcRk1obbbgVgjQ9MpGt2/b6CjcnZuvJlRgghCO4SH
M+/IGLWmiRqVpaRSPgM1kwv/ACUYvBPncTl69KJPKBAge91YfO2TCDKMdt1VYlqM6B9ylsNP0hJ+
jrk9iVZ/Bi+iFt0FhUPw6c/bU2kgDbU2Vl8hZCQfxSXYDR+Y3M3Kys0GbqupJCz6orGzKDHrK5iq
kcALr406kZnp38169CtZsBFyfrpn5wRGBpGdxDYzmALgzPzIyzgUBTP2jqgAQQtp6/qJ3Jz4g7d/
Thqyt1xJnDLtMmHDHR93Hu+YiwHDWjtsBIh1Z9LiKcM5ewXq5sdpGXri/SrhaQhBAFV6HUxfCQWR
p0W9fbW8tbCRWx+CuhA2tAuBAC8BFObkgSk/7xdlNDBD+Kol1RFdecjjDG71BGJDu3ROtEvhENI7
46/F+3oR03db1Krj8x8FmmRxk7TDgjMx5z/y8X1Z7V0wre/Rcxm0G3dhbDVyOiGI6ZZfTEHpnZ8o
1xhtSRgIOme81MgQnojloHKT9W9Cmg5Uhmftb1vZa0xv3+wjNMjzdRCEtDk4q1tD/XPPNiH5jfim
oNJomaXENdZ770oIjvpxE9HymRP2T4Tud/HsZwj1YoodCaHJKJOPfTA8s2nYT+AMkSGPsBWkjqt3
cmrGtCowW+H6c0Vqm9RQgnEky1kTs6lc7G71y2NLTtrvc52FYw6/ftePG3Di7V9PKINw+Dag9Jee
Tg9mSt+jgHW1DYGfcPH/WwjgHM228lDILgVzMaZqjhM245YBNrYeKLF3HGsPFp7bNT0xGE4BE+5T
qTKlZDNWtLFiZjtMIRAXXGFGSieOq2OFR4vvEZruGDR4fMkBzbMFAVWQHw5c9nCjwaBUgCNv6Bdq
fdlT9uIHIMDDGv4behZO93AqrqDB0Ve/kpN45EIGGk4Y6aF3+qm8rkY3dFV24ZVvB8jJoemybwmE
9HPGasa5+WeKP+YLuGbA3g6X25l8wCJVyOXdMyizqK0SK5nkAtZb4MoBK/i7sEGoGP06RwyBzoJx
a7axiHULaarZlvRbjeee7aStK7axSRjf+y2hqNirQaCAGOahJITf/kXp+qnmuAwZ4lrzeCuxSNYN
RV5yurXWFeSqaeasmLR4cz7BH/6Q6K3rX8gh1GsAdpLLjxaqCCir1Iy1W7lmQKRG35mPnKbBTzzR
olcyTYk5MWoAqrT1oWtcRUFuGwusVlBg0HAMBn9X3vJI3RC64lB/2dABBxG9L4U6n2KPD0/GAscS
wAK04xm8QTjMFhZs6qqnEfLzjSewuASyv2mF0FNA0R/cFi9DcRU4el0q9p6ygJrwC002ovFW8JEh
tPt2+McQSK9ILByAull340wTmKBmkK4iwL8Tqco3FVNhr8En9BNSxUQbnjUDGfP/Wi3oKIs4aWaf
4+qmbw0XSb4zw/FTpWhs3yOsVWUql23+gxKQ54+HZLB8F25rAHd3OFbzAOugF/gbwwcoB5lOYb5o
HQL3o1qubPhvuwavKeMyVinmBwoxAxVnhLjHF0APx1U86UY3kE2AGKj7UDeSSjoSWj/qT9hYnz4R
0o34wM2+/Ae5zqJCdNdKm8LEQ+4uEnz90OLIbTsewRwkFCGCntBmr9DHo4MXJFQ+fOBRgBvd/Cmv
XrDiGst1UZaiPD7E06XV93mHbWeuzfqxdXgH8UNQqzRIbDh4nwTujdp1hspxga//YwMhfegC0haY
1V2hYJWv76UM1wABvZKzZbnyPd798dtwjZPbFvleBp977GqiPGEwlTvq23646AHAO1WFfUaIhI4r
Vf8UrbLTr8gwAnx9r43ZPniqdeQf7YXx4rAxsru96HDbDyS06uZPastHgcgi5zrZZZ4C5bsFKzHz
R54g2jX1dxImTt/HtBUlfyoK9wznbrUI1QkijCT8i0flaWRkK7ZRJvwLEKVeUWWDnkVcqjzAtZDQ
yTWpF+xlYJUCcqroETL/PZ9irAvCviPV0yr+HqbiFmJQ4wHGd4RIy76CUZAAZMUZzw08MqQDw/0d
C+fGtLRVrUmtwzcExS9gPvtMK0DRsC/B63T3sXiDEcPVYGLvpjv9Y3a+EClXkUoYf6Jdzm7qNWpE
O+MRUT8OEJrWVdFN8rbWFe7ZEKMJHaXbGFF8bQfyzSP1qz+/7gIvd8qDuELtNzfWX5ndO03JN1V9
YNh53Exi7mSL65zkq7ew6RLU83cxhwEsruRCZKP6/b1kkVH7UiPQOvziYouU2+SC8gc3NcwlsEEx
MrsO0Tnu78nzUVoFqeVsYos4tcNBYxLHB23mPYOyo34m5ibrFBPLSSlXmSItM4ziKESwhwqbmWDq
VBWzPGBRFgcgXWWGuvZinD5GzqkkNYu/7M76q6th8hZ/9j9AEtaGS9j8OnvrB9TaH5pfd2n6eaRY
JUEHDErJ4cs7F1CJU42HDtb40zc5m3KwkXYzgNm5yrX7pPlImfPdtQ17l3sQ+MK3qvM4wLwS3v7G
sdWoHrMf+1WiRJJi5U0jiF3F8inPH4SHoS+ee71tHwD5P2j5aBeoh9yE08IDJiKlpo5/xrkFCz3W
u4Tm9RcJhRd/m5L1P4vcGKKak4r4q0ECagOgfn0+WA94a/5s4l4S6VfXoZHvuImbgUBC7cWwhdl3
xjprhDvtpwEeK1Rgsv9dLL+y8rt8LjWLuLC3Giy2ZqlxsVkcCTZqYk8mxXwl/kYfArq+Swnc5v9Q
8zkf4D2viTgyxvUYCDTdshFBSXLc1s6bVBMtwXbusaEXIhxMahXtiF1eGCfQ+VZ1kD3AFh3Ok1cH
u+7nKyjurz5Wln7NfHqcJ2Spe7mmXBYhUZK2mdnWZDFNcFVPIMwxiSRVPHhUesFw0JfYFrnS5HsZ
Mg9ks++Gx19A0/L9lMTm5J0Y2Omi+lzrqrpVSVNCqbMmlekTX/JCcMwYzFd3I2CVgMMwdYlDOBF2
eF021otTaYkw149SMH75slA9UjitlHDlfTghya8+SexvVUn9AeQqg0euUKkbugI+tokVJ8gKCBqg
8ZmXB5u84iyp4ECW5qEbHbOKnalR7jI/ET2iiC+zM3ukAn+w5cvUPHL25Zw+SsZH4+nM2iuN3oJf
1g1jmeyRpVoo/UfwKb5Ng0+6t83ogAccfRmxx1fUo4djK63p0SG/5CoN2ZmVf6RrkZV9VowCT/2i
VWfnracizQlA71wLwI4OAkhhctzjiYK2GflbXEdNnjJah3kKtQGL3zXG7sJatpfaMNCLtcywPoiy
UFVwz1yMIgnim94xaUdCJDg28PO48QvxWI7QD4ZI3EBUmQbnHC4yIJT31GISShE3QmXo3KiVklSd
pePDri6CCwpqqc2QpN417qqUqIA6fN4quCiZPv9YJPlrP0Sy3Ol1mh3FPdlTtpwxHJMWldn7vaIA
/HcYGPrRbCiRcV9uLKI86LO+7UXZUix0Yp7FBeYBalMke7/WJRKLxGFGpiWUNCIcqIcG31VQOPRt
sy6aZ+Cq3yQQHgEKOcHOUcyC+x7Nch3CNik5BM2czotZA1DAqVpiCgbcGNzeVLF8Pi7rbJfHnbz/
FC6rHQ4EKENTkdRCwSi3JSTmOKhgNVg7z1jZtjQFI1JZul4Gx0aVo1M04gcP7yY1BxO3HD//r+Vp
o1MHL6wg7+bABHg7ishCjQGXtG262i++y+XVSjKW9AbFCQtoQu987IVJ+6rCcelC8bovzRo0dELl
/S4NrKxVfSl+e8b4Uv96nhTVERFnkxDBnFYMAYZuFOqlvFGTY01BhuHDRFuC3nthEca5Hy2LI6Hv
fXgijzQGWfrTSXeTT0FaRU+5GMozyDfF43J4uskPohhrDP7XAjtbBbya+mypJux2QeW4A+SoBcUx
ka6bNqEoadRef0RJnBM6Ym8EoM1MXsLosSHmeAkhqiCxsjvYOi9v1381l4Ly0KS/rbohTfW5NQQ9
1BRXbVnHuTR7M0f5PoXSOt23NyuOF+h0Qhb9tfHkaxviPcUH9jHkzclDUkjidZKFgaWC6dJo90lg
JAa+WVidP2z9yNIOXEfWD7LGDkQSuO1T9aTFASkAht21sQQPeK2MKskigmDO2NLEtHkP3ENQs1MX
oQ52w51DVd4taNs4ymCY9tx8Q6pGCToHGNVQUkmars+weh2QB+4WZ01bbgPBU49R4aetmi8TBJwp
PqLVXlpTWcd7+OMga5Ah7Z1GahwaXVPDCFw/2Hffs3VjlBXX+bSR6Ly6OapYdS0B0TAErj1OqUEI
uwaaBeyxrYOfGjas7mxddBl37ZgZUH1eO1jkWPG36Tjv8fXLKB3jaLaZCZTiHKSEf5WtO/KK7G5x
cLO2BWsXqIn3jAj/lPFkpx6+5oEpJM7HD6Q3+XojfvIMp8xnBYIjlCUUT8pB4DKSVvDVFPNazv0O
5aKbyul/KwhOUqkvIscrwhdHkY+z8Wbs5x/8/UYhP/Y3fVMhCEVyAUI+5c3s4aJItHfLL2kdlhaw
Vi7PNXB36945xGE+9oVv58rDeG8V6izBe8q2x8+EFuPyeyiTXEoNUULwCcrZ/7sWWnfhkA7q3mh4
ZhKTl88O8SjkgMqW5Lupm85S+jk2Rt9KvjcIETBHFno0mbCKSwD0ObrpC5g8O5o47mx0JRom/xg3
X+/M/FA6WbIgzRuWuI/VL2PqnA9iV25s/TY81MX70zs2jLRfpk+TpLk/IRndzBdKcjYyKY+PB3+I
Pm+tMrK5LbiNkSLcd9EUULYy/y5DXwPsTwSoM/cNnOB0ZKvx2XBTeZPwLXlu6rjuzumcLDf25n0j
jjzCf1fzSQDO31vImYGtjnOd0s0cVO4zibWIHvvRjjGFqoWu/U7XoPKrWLOu9cNK6NGDSgrHchVe
5Dr6LNiQ3qHw8/XFQU6zdHdJ7KkF+IvqD5+WYDWEzNdtH/alElNCyyVvohHRfN7DpLSq46vT0J2/
91VBArSvyPEjzaqsZScrVBffiNNYSToGzbLUT0Ard4s+tUDRANy4ScUUWO5617xAyyG7SnFKaw0z
G3EKAWY6+IsSnMzEr2qYuxaumwCCJ4vkHQbPR7DclkgXlsPRN8DgAae6Z7aZrrmv6Ssjsdl/w6JI
Rus17vMeu4Yr1sjkpvd5WN/ViZ6/pXhMNwgrsv4IaMUrn8oe0QW9GHBGffQNoTGT2e1W3dHThh/q
vq9F0ZcupwfP8jYeYrtgpjSnbwGNLUcVMbXv0IjznUGdLbPXYxSI/h81qph52/Mx21HycueQvh9A
pnw4eIf9rd47jo4bdHrh950gthroKzSZvCeANOYpzWrRueueAFJeI5ceRFaeHibbvS95m3dJSu3G
3FkIxr7HQWQXOyv3cjDOYFvOJcOdWLTaYgNTTPNLrbgLv/svXweklxbRm+Mc0NBzA+m13zovKBp8
Ksoi3cT9PmHof65jtoP9ycZwUba8qznkIblzQ7JqhCeL6d/5U7ksoOIhoqm39LYQx02iHd/vuiCn
FGxSP3faM6hxZh6ssvHhNIRWeWgD4bQH/PveD47PFhidbqJZFXfqNyj2VYHiLKN/VIiqZcVtkF5Y
8FVwVwCV6eFX4wA+CeDCR3SBeuS/4R8Now5yUTQa1zT4AuZ6FGkJG8PkhhTRGlLBRptG9cOmIWoI
T/zTnqL5psrMehZOqxtQvnCBed/pctNcwXv0L9g573ebFBCP9qFanQGvRvvaPN9ujywwglirN7Tc
y8fJ59uucgTrT5ai0Y0FT+NJdWqD5tpvW1Kyk9EuDKLbHIbigy4BUpgSncpb60uqFQTR9S9o7EoS
Yp+xGe/Rsx6kZ832N+Nmk3tjJHXWoAZA0XZtmVQ+8RlfZx/e7komJhegQn57rJA6kHCqOn4t3Oox
03ZVDuU7APN4ycC3255d8YqQywbHXx8cAJxRrOq/056UnXIxONPwJruSbAq43Sy593wOZZcdloFH
ez0MftBTZFWJL4D/qgeXmtpethAaU5DlB1jOqn+J6KcRxmckGGHfmMsB/I5TRuvOpYyMCaXmwVCG
1bzmUX6IUD9g1MzhKzUsdFfR3knItdWTAVtc79U7R+Wt8jMORxKRnl/t0nSWwhbfbY8LV9uM7tb4
S6C83Mex28uGsGpIXMeN3TQdFBijfZ2poDA9I+jJgOJ15Cs1OHsneSIKsnQCf+6XA8NPxJEqQfKi
xk2fzjTh65QNlcbMCjKQ+QX8SRZw7Mh0VVSNNwgR7gre04Xwabtx4MvRMuRrgXMoMtN0NGga3CkK
L/8SS2XtZcekk6fPSVu4E97cy7tUXoFMqZW2YwlHptyR8lkDF+M0owcTILxgfXMQGbQg1EgOulxz
h3JCY0KGLXWKtbFUWzC8vEwG1swp0II3UfIUq2Y9IswvD/40t3QPHtvNNlT2DWb1gvUOns/cfWqI
iQU3gXqu1rKc7AAe+euQbczKfwaMaGrZoKKdRhT7rddwgrVFZvKs6m4K1upSbk9NQ6Wm4pkoB05P
2FJoVVFL0w41DWKygTaGuDf3A7JpIL8wU+T2ktMI4wrwo7L/p0IMVOMxE/zDDGnLoeICWBGcbZea
YfL0ZSab8eIaaSvMwEQukn3JxHJTUUBX6c0XEv80sRIzKYL24T8r7z1fCapOiHkw8ZmkV6g6aYTz
ofzHRbJoweUGCJKr5dmR328LNjvoXoa+4804FLQXC2Ejo/PBE1lj9Sar4ZHZo6UJzhC7q++DYkSu
EWVXndazfDmOMZGrVlTi1kKxAvtQm9FSVQMK979BH2WmdZiK69SFghFrJrB0FdlwHD4llamrn6FQ
Npr2LLg9fYVEoPFWt7Jb/X4enJAdhwbZcg7UAjrUeFsmfMGRh7T5m5MROzkJmYRE/YxMOBpq/+Ev
/fLXGpUJOaOM1XYHISmBSbOyEHjYG3jmxB6eP/0Rt4NTdICzC4+KNEcqKM+1H+Evs+ASOm2m2xJQ
Zf8D8R1Q8Rv3vk+gU0XG5FV7k5l4nLAK+xv1sGW4alWZljsW8+iat00LVoGUNjyAS6uYWwyYjl6b
c0xIiJWkbrYaEIbb8D0mDZlpWPd39xmPztdmF+0V4wN0mxCaydc79HR254b8mMkfcucOzMq/H7v3
9gasEm7vEOSvqMNb0Uqo+5bjaa7CwcdLwCEwdMMnK1Ah/sJQsHIzGCuYhTBanK3uPXOPN3/hQVyR
y6Zr79HhCwTd0iY9EZ/GCI96M1MCWYuYOmYRHRLvuGTy5+em/vspHc6PV7sQkHvTgBxIEOx0/2YJ
UNpGlmSyuL74nqwnGkKECTqfD3xWP9jgXRp+aD0W+gpbJ3WernTTr3u0QkWWZg5nCI7L3/Z+fN+s
AGCz3vDfR+fRHDkLX+rc0MIM2ocSv5z9rDnmkTnwKou28JlvcBHP0PzRlwYKS5s9HplKHXNM/gzp
8o+aAViT/XGxrqqaNohxkepWc4EdHyUVjBI/pkfXPTF6vpFjZUY6wtQuGNhAoObXYxBsJ4FdhHJU
rBZt4y8IKq0qhKZPV4XIGvkVFC+CrHih9en41SaVLdQ++pohT1WzuYgB0rKS4IXTM61dep3vJdzO
1LpvPt9FUN1uxGzFW8KFuiLa+5w/Rmf6TZPf2LjCXOY6rQMD8VG1+UNL5jOYJe7v91wi63MRmWqe
r4EBpsUd0xIkDlXmLzVaJMHogn1upxnJKzSLKKcxjuwNdEqXDrHyH5cU3L6QXDBtuJJSbceXpzIn
Piq+fVj1rFg3NWPm+heECRaQ0Sl3O3PRlkT4cMxxa+4EVldnNJNn8HOR+MMp0CXP+jLzEYBNwE9E
MD/zke+YTjD2E9w8Sm4oVBBw6aJ/WdqY1gRkuF8F62wZbOL0AfiPWx+pvIiSujfyul85lUKs6RT6
EpjorYg9pB4Hp6D7LyjyZxnYDE9AEe3ZSrUSjCm8KdYMC9Rn4FMpgpRYe90ruoLqAwbAO7xuUkWi
TLvzqedbJi1Q3dD6zo9oBI2jsulXNFnUJcx/VAVrox4ShMFvXyQW8eHPMM3qOOMugLoIEgh8odTH
beNyQSpee/6EZtjgUs9y8wCvnKTEHtb3lVpkoXNlTjzbGPTfbS+cBgNltiExBqeDQFlzB9FQBBI0
njVU6Qg8KE03oOS0sx5gjwLp+9h57vFatno0EI4GW5MWT9S3s3466NS7dW25e0eAhO4oNQSwKi1m
mOW5lDmndxWOW7nCuqxSLU1C+TgA75FkeW04Xt5nU7g0cZnjLaITA1Xy7nkxg1AlOlss9EqL2Io2
NO9kyrQILRpAGmrzDafeYLI9ENhkWvAQLrQAwTuxfawFgOWIQz4WATqm0TxF8SREbHCrMCFSvbJM
K4Rul3sY3HWDrav7dH0I02xbIxkj/L8VfciyVpqMzBW3ki0IEH4+QP1paGGnBv3bUyfdPEqOwADx
CQuYWAwzIHWiTgkD8uF1qce/E50vpG5oQrZGAv1HXaqD7D6SVjTnFgIObfPL1CtqGrHb1rvq3wF2
S8smoLFToxuqxtIPY7da9bl87bG24N4knDHh/iMUeJV1j60c4BWVwzsTXVYtBulkU4btDtK1CPYf
JAh1LLAT1ioddP/lvzbOWGPfkzIW1lu6i7gXdTfMSrw6wpx/QcE89kqpK0sEEBns/N3bC1JsWY4w
DsdbM6D29CUD9HgHhBuk0jE/etCByAHz2Ass/St8pyahkA5b3k3AliEMht7afmLSDEpwwdjE7rW/
AGah0Ohs++A2ZWi/a1yQ7AWpWWy6hQKWbT9a9LTwt5XQiQVtjkjq0ezd3p1Tdts1C7EWxkP/uU1d
jpAS1TUhLMk+9PHniIMyIx3XhF6sgQMBwCK5DBNPQo/ICP+RZhCJZUWTcWWG5nsUOrjdiYnP7MFX
dfbflwBF88oqOy75dUvYmcXpN+TozISb3PUA6C3zNwBQgF5gTeD3SHRtLa8wCqYmD4rFlvhszxe2
jiz7iyVoxWSZPvyYlAJ0cAQXe7v2tlv8F1mUvVVOTyTuh+67mo0FK4nU77DXpIpy190e2RmfMi2X
+jnFxbMwprPYLRpPnXwemyS80mF4Zn0cIUwqFZabPSVKZE0a3HMTgxPY5Q/Za9GrhR1O+J8JNq5j
QmAbRZ9rwLgPh5LayHdFsS2CCkJJMHnO4nulP7CMz+Xi+DotrCIa6xgn6icEmqRHWEeCPyAtQlAJ
j4m+udjvgOsHNV6lL4wx9PGJhIFqvmsZuAalFXCprHT8d8j3f4DsCE61pzkJscH5IvEMhzpkZO3U
wOe3IReQqn6Hy4U/jyZ+0u2Dha5YsB6gt9ksFIyBcfFmBCllzKC9MHE9Yv11CQLXkIMF8tuAOJLq
VVh6hohnbbOu6aMxTQ4ddDoM95dICB3Oe4hP+EnjcI7x2ulqO73GBzq1Isrlyv51ExyEd5g12Iqx
slyUHp0HcCbXXZi6W88G2t+L+8gu62Kcomv1QVTvUURCStAE2Vx7/AeGcOdLJxbksmAksJYrEQF8
vh5mFNh5WEmITVf3727fsElWLw8g2rmK6+AKSOzyq/mxX+PPxjaqHZwXP9NtJ0KTdOV5lSSEkTMh
PXRKdPGRQNsZybSNRR12yU/H3KmwxYdGVrJgP1HqAqno0Nf2R1/chPQ3Cw4bBcHxqGO2WySDz0VJ
uijty0eUjogAALA2BpDi/WzybuE/Rpn4E8vyE/3vC5yFdSYjPEaZUkNdZJlXiRvaojrkWMqef16g
OmQz78g6LeLi6G7iEV7LpMQe0zKNYrldmJtn1d5FtRM2MUtdqxW3CTyEua3fsMJ8OB8nYQv33ky3
xKyfISqzT2kHg/YGfdzd1whqXkoKa7R6TjYCqJ8T6t3FqW91hvJnwVyiVwrulQqqMF8XacWnfadF
tb8TjC5xEUch8fAH7Prn0qXvFMTS1VjK0tHJTM7Um0ZbhxAtgkaRXWGzFtueF8ZVYLWy9cEfsG+F
3jlUm/HiIdoyRS6EdtMWYKKA+zU7FVsD0D6IRztRSVZYy35M+5ft3YlyzxGCVeTB2k2IuIe5qQpJ
b7ZRvC52wBhDemZzltpemq6YrodbJIguHI3cqM9PebANMFTHOaoSRZAZEaNou+2Z6uD4PmabC97x
JUT904Rzn0vRjpgtth79rNfVKz+Jwe9G9FQR4V+6VeGn9HsLoM7nwif3F/+ylPYN/DnC+nfg3Ky/
dQrffTcl8p1KSKik6+B/p+od68eGMNvSv5j+e4tY62SSzxUqrO0v0WUbALoWTjAsgfl5NeUISVSX
Oiz0TmPp7+coKBHcNaZ3Rg9wI+KxGnDVfjEhEM/pFdGIC2RiyXcRKY7k/NlePn5AvIXZz0Cregx6
pOqD5xsNHy+Tt9QLA5GA1w8VHp+2yvyF8y/dMuR+c5Hkzxuow+ERxv1+lfE1poVsRbAdTdt6ySbO
cX6wFI7o7xxNgfdWTjHKGELTs2jo0E2Pp+aJ7GKm0u1T1TIYp4h5xEAwmdD601zZWcDoTIU4nboH
zDdMOLQLoLxApqvHwQv7mgDxGWPjB2jGGsDN7G5ncnTjA59yupxuVgHkYfEOLVB+tzg+ppXOSueh
jLN/sCZedAXTvx8LL8ffHwdlfE5alwVEBBjSjlQuDPXsw7pTc0Xrquqm86QcYge3g3d8cXXf5IzF
C9Rd0vEz4HnVwn951Q7nl9ILs0o95z2EPeERpWukSziD/5o4ECe7GCCGVCTS8a/57Vw1yNxkQAut
mnPOvLjM7cLrVyEwD4lh6jRvD9JaHchZAbEpB898/38VSFmk79b27rh8tVkWRObaDu8ozobWdZIL
vE1TDv5Sf1LoYRi9fZP4PaBmI/qZoJAQaiwjQuYinWazqQkDN0aPEOX5xMELMfJo27C+K/V3wn1a
PiEdds6KY2wdTsBDvhvVYMpr4BH73G0Y3LaffL2MJN33fCrBNhx2tZyiZ18T+e3/3Sa6hBSMlyCM
QUZORCspmwuch0Io7ei4WaAsiQXCJZ35sdDNc82hXc0EoR66ba30oQBjdih4QiWRgz19pFT5drEC
nIAE0Prsc2iOg5vAJHG0oKtj5GeFsDQ3rEQJSSBnJIFJ4ochcA0W4EVzd35OAKpFRNZt2KSDR4iA
Ctb5eonuqV/EADCm71ORA1blMSkmvumaT2kvvlz6o9WoCxgTaZMck1VGpzteQvXnWlHA6LWlgEte
dQp3f+ZH7HzQ0+FIcb6D6ASdwAm1E7SBwZJcZ4OjWt967majWc39ZbCHEs5sokgSxcWUHESUz3vS
Tm/dk0uXtnwNlPw5nLF/jq40xqf40mUsUgT5vPd4zK+2Mu/eFsjRtuiyPjZayFfdRwiGS7Y9xc6E
DACAxh8qGCpLB/oxNmaDT0FREgKxtOg6Nlem4Y8aKK4VAvKlv/yCd+Cp5lqKTJekXDYjN0iPkdgp
mw94JPj0jS+xFC63ne450Nn0gcKTewXH4Zj/i07RExcag8Viblfs52YeWp6YdsgxtAhp6Xaqe05+
9QB8OGQ4dW+EOyoOEPh5UW0tSCXqbAIZ/qRLORcBYAgA/8cuEPSrSUmNIQpu8Gmm0jnMkNyHR2f6
wGWaqgcmxYCrIEb9xyRr4y4NAPCqjikjln6OpIpHv9Uveky1jjf7iioXFQQxtfiAczJGGc6FAaV3
TxNrCK/NRB3akeZb+h38JXUdphaIkEm6vO3IxCmokG9wjKDLQKgfXOHIoii6InvVesMT64aPazll
7huZSLUexhKLzYrfdjyDaS7drRIig8qcseBCaJO9c9HQB4wMjeoqWLQLOqzH+lzhPYiphXOO5BBp
PEjdZyOMkqrPtE+QgxoaeQ6kooDs1X4Z6zds4OoFFmKRHjmR+c5W3etTMmqshtSHtMZFkNsyDnvL
RGSwYJkSP5kBk0jD/qknu7IjxfNgZbsRg8Lalwzl6aB9ICPNG3im3uN2+9FebE/zRBvJEvr05J38
qpkknZJb3otWlth0ANjHUmGkjCPr+4irI83Z3Rf0QTwmUOyf52fFtfNgL0zkZmEKNmzoBCxy26GF
AW8Eh7vqG+REgOk2K7AyqiPIPE5yRgB0rf+Ac5N9B5Th1F9C8o0DhA+tpKDTsljL/5UxnK+bviem
q+RZj0h6u+0I4jMQCwHxa9AafoEzsaNlqzhBMWM+mMA1zudsHjxMa2+dYdXpgFKc8Hru1EngUdzu
yQc2YVbzNSTQJDoib5gRzNYEJKI9Y9hF0zp+cZvvYPGyl7hgVGowFZngzAV9tfBclNQ72ylsciZu
RMV3w3SuAod3e+8P7XukGWElaMAVGjOpvhWB0MHT6PLiVgrww6tFJVJkRNuu/4f6sxMOm1rgyASx
TrkWIkm4n+lCHc2n45pxlxM/GuvvBkBH5H2j5/26L0gXOYNMK3BGoSD55CEE1VB4DqZmc8CWE7kp
3/Ag1tq8LgIu5Bb9hYW3ZM5M7GLpjlzxpZlTqsRT2lhmkWw6XMuSAQ5xYP6AWkYP4Ujfj6R6fC+8
k0DS7/YdJhngRz6EDFD0oWdqaET38a36aYg989RdG52241XSp+Ikn148SoD+BIIJWrjVTQPwUVfs
/9+TSC5N640AvOI71d5Tm4Ib/tcH9tTZ/iJf+oo4SI5apH+C67RWuz+/29WxKr9279pqVOwJMhDN
CwFzFnwb3QaxnyQMOtIodAyrRz56z3LARto4OciOZvnEpCCyxfyW8/q4JxxznNehYMwJDrbeNM7O
Ln76tdjOfO07oc4axzqO0S0go+EuvR6de5Czn+CnnWlZtkmAVWfL/Jh49gkmIrtVIigzaxL+ANoj
PZm/sKB2k6lEPJ4oMZePewKxpcAQ5cx0cIKtj9l9YS+pAs8YJ3cvhrWp9PI1cqw3PrUrZ16mGU9q
kZSQBM8VN4xJq5XdpbDUPXFxzkGQ5uXc1I9XkPHFbPBTC4p1pTAE93TtvIrf8Gzpqb6NV5fx0VJZ
IoZtvT3rzw191ZL+EUe0Q0BsVv4BXryV9oRFqu9tMtPiFF1FR1/tpVR4ylZ79Cdfng01TExXZD3W
BAA7BGkX42MKDy4OCrRKKnQeeCOZUWm79Ts8SMCjK2uEhaBQf0BPPFPC7V0cSlKuKJfUp7+dZZrG
hClh7zfcvMpOPxMlxml0Uh4uhMQceu590GUd7/9X/FP7E2XPCuTEtAhdTcNqgBvIGfVLsJ/VD47l
Q7aCn5asYSGCO63RSZ1SRsqtB5wuWp3UwWp60PVE1J6T2534oz9irjxHUAn+sTBzxqLJgDyI/7RY
DxKtmtWmJhtc+m0g40+RXKSC0ZW+aXaOsdxz89xzdkX394PtYRJtCjaOMeygFGAOajXDsxacfLtF
ARMywhZGalY/4Zw0uwQT42LCE9GNvYjTQRMmrzI3IngrvrIFv2mxuohhQa2mCAHMQsYwLg/18s/K
vwLr6FXWU3PU2wUbAuKFKJpW+5Ey/AwTP9hDvTHt/vHSpP0J/v7kO6VlZZQovRskvo57V05EWm+Q
Bu/Ebpi8Ocv42pH++W/saPfJ93WryUirKgO8zoyQ/2G91GILwZBEpHY0TxtDbZhIW0qHx9l7GJi/
KLRVgWBPeNxC+3dExcHpxNWQkoxhZZeAART3pAphpyagrdtFHLnx68W7IX7X5941GU1IpUUHtacR
+Mf+U26l5rcT4xAzwOHRbqqz96yCYX8xAKeS0+438WHxQ3Iy8muBNManJYhlc4+uQW+Sw/4Jv3cV
7y3Nq+K6CWBbhltR1Ko+XPICmwC/cVv1NYpZAHxWMrmof4N4dUfXkATnXZ8y74FNHCLlSmWdkdwG
Qbd3IeeB4zYbYo7NpWwWDmJWTpc1tuE4f2+C4IsQFnYU4g9CgloK+P5WJ9SUYlZI1KUkc3NQaiVQ
3aR0WjDYfuCLcHZYt7n4RE7DPIJMuDAcbVMnLB5IFD54FTN9ARhYa1bkZEh96NGarYyemfvgNkcI
h2Q3YvKxILorEWyrsjDPrvcvMRlhqe/zHKsJ24fzgSkyV1gzm5kYSvhuL5/o5ZilxPfYxcrlgNQ9
FuCBpqye6sk3yb9SWb6vef7HNM5l0SS9im8XIKxSwbwfgHKnVEMVoFz4fG6rM3VkoaJAqTiUInZg
yi2TtJO/CYFMj23dOLWSgij/6oAM5cbE287r5/6u9LKmYoMSMw8EBRFuTsEMdowhyoOu5OC7hkmw
S3pq4yzGveHhyST60MfIsyW6anpi/VQylXEPzYcMk5U3/hPKGSLwQ0h/ei3Pfr2F6aMUssOdGH4v
N2HwZgCP6wRzuQ/pCHdaBjsN9HKE9nQoa39Rtz+5B6NVa9Sb5RK3i7Asw8WkjC+0VHSefdMBdTsS
OijMu1OEwEYu0QXrloNCskbcXQuxGAvgsVbsmtuyYsybgabDGY+2MO1NOL4LGdvem4ACp/EDUxYp
5cwStqfHdeyZiL2zcstJOdT8cmDBuF1iP1FA0X9ER+kCouAdBjuNXiNaH+RwpiVByvh9z8gt3mCH
14pMhHyhkKdCq2DGb2IXJyNOhbcCxIysLjcGqx6CwMifArg1hYLu9w7w5dGSxB0Ssnu0kb0XolyG
mtUPFRfC4MmaEf6r20Ai8t+0q6rHGuJ6eLM1UQtwObvFisiUApSEHCAI3Q9lZ+ZOYOdGCQH6NQlV
5AK6Xb6cWoDfcopje/hSTy5+kZQYhkg+TSEXJmZOLSoMjgKpdkgVm/ojOV5YcR+rSbTOOLm0rEtn
HpiOQZg38CO2bqbiD6YYk8qBas96gveZrkrCai53k40oovvaE48dKZ4tqo7tulyy4ONBSoWUWxCx
1MNxAlgzPmd7a/f0NVU8p9YvRDpq0MT1t/z7GStsMqvW5uqulVx1b2WbavO8EsRpFMP145cROxVX
YhUZNqg64lk9PwdrTSnLav1ZMBVWgCh0bm9dv0vIum4mX65RJ9OWWMaN5zF6UKvpIqwxu/4Rmlx/
Kl7+NM8qqfHGGTD28rlKa8PdtKZ2rHB9pmOhe0OLV9JwUK2ps5hGYYgsWm6floXp4LBotEzfhZ/X
gc5YvzZS5q8lamAMIbX1+Gg5cuVRV2Fv60sPEFzPBNL/CfXV3mslPHHt2UcmzQPSrBzVvGWKhyhl
UQ1dwEZcOjdSfWHNMMZmOxshoHGnKdPxCkr6fjsbe0HrGGeJF6T6gIWtVbeF1xumYH7evV1nkOD9
fvL3c2U5G1NfAe20mSaZQlBgw4BnUXRzSpjUQQKi26BYsUrqz8028rRFRqxTuE7RaYmNFz6O9M6S
UEKYQuBscSc5E1M/l2DOv9ntyqW5Mqb2AbfmNECfiUrrsuL/CiNdFf6u0XMOhThsZZgl5IICqerT
o7iupyj0IdOJZ4KpgEUoB9Z6pegPymTMXcWEZrGLTU4iV7X3kzH59N0Lj118pcTSsXMCiqcog3q7
/nZsNDCbKrPqr/cLrseE0WhC6yrNH2htozJtTkqnjEjmDF6w+i4+42Kf+uCc5up0JHkC7Q+WIj02
5fzdN8Czo7aECkehQ3P6lB+Cj4q6mhmR/WdcJ8Wzh6mPmUz4baDE/iwksusq/9UD71yAqv6HHO7Z
I21dSkQsVyH53bed6pzE3cetoURlWjCIATWJ4+khYqSjBlWENNHUlPexWlmVEIp3vUQVeVUOsPxz
uRpZKzACEmU9BijF46urrwbzKZI9LEpmDT+P8nPi6/yAkT3fGks76dPoXdGxQlK6EUphnyrymCfh
FEsOfbCAezi0AH6xX4VCswuQx0qoH9t765TzBwLAyphJsmiJACZvOv3Y915HnCcbiLpj0SZoUeWX
R3V6UDqvgTaECg+W7Plu4ECm+MVD0aSwBYwaHEBwxe+r0OwFBREj41Z2p2EI/+X8JMUqbP/aB8b9
WW/dTgrZIR8bIvuh/0tQRQD0ZpXfa2S2d0dm6ZriPZN3cQpHNSyFGCpCs/AOXTBn9sxcjPEKyUJ/
JtjMQPIL8/QUj6Zd6AtfyS6AlHT2O5mCbnsIPz2hvqWVOz3LqTLYxmePoAIW3QFOm3jQ7IHnxkWk
JZCvgYjPa72c51OErHLopUnNaW4Px6inT1JoxuBGP9G4AQkPskS/1zQ1l1UZ1evrMy1nDeBp02aB
Be4U1mWWWxwVDxCGowMnJuFLRFD2nK7WL4967vY4bNOk9lmjmT1WsBQbWXN5W5rXZ396DBa1vWa4
LbkZcKYFgCU+XTHmlSshT0gl6BF2nQQgOC7J/GCfdsbVzpMHrnoc5qMARkv67Kr491gDTGQLIHzS
2cs3DQt5qmKbwpw+16sk+HYELG8vPoZZo8UgfJoOPurMq/ffHK5GMqIHgCwB3Ej1T9zsHxQf+3FB
/qB3uClKbd4liDdtpBP0vg5aUs1s0FqyRZ2dNk5OZWQ9UKIDw7QFKtig5SUswomZ9OGlTk5rryLb
JuJllM/tfvBeq6FZAR1MHQbKl/q/Eh1X0dVXelcyXh657p2I+lAtTBOnxlNQTczqCXosta3tGIwz
xMUyF1eGQRk3L+jYj3gjSkvoERAIQvFxTtenJJu8qn/qriYVmjqO2zFpg3U0qHORORxcnntpyxZS
DscDDPyZiKBkcuwwubz7m8FAueAbPHjobgH7iUbK6II0hA80KA5La/UfnuOjFH1m2Y47a/Smoe0g
g/BeV0zmI7qsB5SWbBtdcERxWXJxQ3RWk1ldpOa/id1N/o1ET16oF3ikV51ss6aTgEQpTmhmDwQU
q6U2RLBKXZS7oILv5bymDPKr/+hqq4LYL6cGvRvpB5MUXIbzc/5CihTRMQ/++9q+JlrC+4mx9o5a
kc+m8bBS8j31mb+Z76NpzzjNP3Y2PCZKy3nI72ZcgxcUeguS+UPl1pMjh6ViJw7F7GS3DkZnQgu+
u7Py3Q55D4i3/U3fYOzOR5sdg9B8F5xAhzgAnYH+OuX5+goaUWq8M6eVFVjU6RfPSvZqEfKbfNhW
iml6e0wB02S4qZcx96e1DZGLlf7FXsNGyeBL0cgUdML/M9hUHJVBFHk4BAv0sCPyP5TKlvOGuVf7
7ziioMh7OZpmxnfLeTIokX8260+tTknolCVWUev+S43t/Mgld5juAopCY9ENx0Cr3nMOAiYywDqJ
PAQrQYdAJEcBud1lCVDRHtM9ZuWVJqNvI73O6ehOkkINy+jQ5dh5ZOmSiQPxrg48rGWxHBXpfabc
xDUVw/uJFRJOaHaBvXvAJKBGu1AsaDhApUw8o9c1jmAxyhq2Ve2cvkpwOTUZM34+J9Hx6M3POnt/
eCwzhL+Mgj6hYbsFUbWCsR4KYIvLW8HDIv3ZF9/Fph5bJGpotVXOpHQB+UNfPpsJJix0wR2MEH0X
KSlb3P/XFWWZ1/cRl6ZL20SsbpdlJjUz4LEgVCdJpzVGpwTo5x9GTmibU8WL1jfDsLBrEn5lfZS/
aKdzYkZqi+snqrcVodUCfk5+Hy1WH/u6fmgtTjNg4L1m5KmCNhRQ9A5I3nu1EtfjgqQiBRJTYE60
r7sBTjtdc8vrmL+ShFEsv2r/ahlRRWIdn+Qt8TzUu2CRn8qN6+g3JLVxhc0VU6ydld/nP5aYPqhG
mgZQcgSduFUtAAveMO+dtWYltn2D6n1QbgxS561o8rpe3YhgyQX8etR+2lhDO4GHTWQkfa7z9y+p
o3v2f3xTEhbZs8ZEkT6WDni2QrcWkrEF4lZwdRZtbso/DSrBQHlpfnMg97PyU10dpbx5vOUYX88i
nijz93xz1KwmhzraXrOKJjxPOKXSw1bKWKuVdm2N8BLKXimerbVoOs2+iarCwJjAEh57jG74bSXY
1B4PzAS4kL1Vhe6U8XaOmBqAfmQKJOWNgZQ0yvGB1FUiPE2TLyIWDfQfpmwG6xMeyVAFyevKaW66
gLw6XdNLjDDIh7D+kQP87h37gvlaHgEIHigZRoX68dIxbEADn3f21AhsXUa7epDfEmsSgksKl7CE
yiaMGznjjmDxpAJsd+ORAzmvW6jZ7baTYICPzx9+TvbnTqXV/KL+rcxQZBQIxL2oREVT9N74YLjl
UeaWCTK8QYdET9qC6fVphTVFtJ4VspqZ2OaGixLjx73Q/26eujByyPK1RfwcJe9KjQr+CUd/tNYg
nA38uvKBUU6q2maZHVfsz6jz53MEkfoBJUgSVoylVDdwvJZ1eZxp2XXGnKh8GLz3+8Qcbc+xAsMX
li/KL/XBewPVSLZ3jE6kaFdd4ywrzWnWEZKi0fBQqUXTpIvYPrNV0CmjC279ouciTt+NGCnn4o7X
sT760IuCAgSbbnNyCItAY2TGdwhNJYg9RQnmmfOrPYanBg6D8aEw5ewWn5hM6/vm3omFPwc+AiKX
eYV4qqdTUGd5wdioTwK+27NYUs8K71Qm6Ir1OnyQNitXiFpCBcQJmxEWn0r1flrvJeAnLBB7bcnK
nHoU02jWfrlFdGo95YnGmAe5CgCQfxx/sNoTPhDTP8rlx+M77kUxYZ1TqRYfb+BqhgqOv8st2kPa
8thptuVBRHEy+Ea485t3mmGNHOAtfqGNwxBuc4YwImdJvL9rm8VA1zUjp+h7vpMEGBvOtLF7Yfw3
g3uniS/CS9nsqRfw5Epzt0XrBXpAIeM32pNAA3vFlvyHhwfASH99R7LSLsHivw79LiCzNUdaRzoq
KbYDSPrAfPT0tL96Fs+8efJK4UZKjj1/CTaHCstUZvlibJdo8akafvfGZDW/SvK+91kfM6IwJi3Q
ictpQEWJbZv68ZDcmRFd5Inj61Rt0LtGdhB464CVo5JbcNn2wxCOveaCc7znI+Ae42jcz5HFNXI6
C9X4Prthnl9sqPLf3sbSewGoMqPMq68rLZVr82nDiwpn2e+v/jSK2bJYi8xEV/Dh4nQvCwxMyw2w
lZ6EKgqUG84SgpQQVbA1kGP6OyzaOq8oLzjY+sqQVg+MKTrR4yrA5UF3eiwv9Mxp9Sa/FX/p6tL1
7QX5Qi8PaYLPr01wczZlG9hU/GsUuWFYWNGIOgqjJ1hKvnOq/tda+Ic9dLLVtY3PqQt+l6GhZmRT
i1J7wDi7XXeo1IOY7K+15mQ5OS+FungzvMdPhL21hQdxVtPUKeHHSBj5GyPa6WKRIwVZYKKi58HJ
FD0Q4QXO4FCMJHjd/HnXWnqBpzdsG2+WVbc4Orp9j6Vk/64nv2jGtxeRRra747EFDGjgXFcoR9Xr
ELUMcletossyUAC5RNNsS8E6rdp4IRYfi0z9c/hwQoqLO/W6JfV1YoLTUcDPkLOvpRSG0wG12clP
FI3bnxpUJPV7LNPTh3ArRrtvYs5oOZ1FhvAJhV0PAn3FQoecB3oF0pjbBPGyOQ8ypMB+A8iNMcnX
EI7jVB2gJWv5uutqoWBa1Nr+vWdNPyO6nAmGx+tVleD2FpLA0m0CefvYZC8V0mNvFP0ZLvBjVsHU
zfLpMGyt7jzYKnxZv3079dOryeiWHZL+8khqn6g3NqGMvf72W0LSKvgxrTI90+3u+Szz92iO9wn4
E/GtYTpye/f0OOke6Q3wMm3K3cSj26tVVg7XrNTGi/qdsKoNkpRgnshyYuMvMSQCETkAn/fu8/5f
EfcgllRvcJEP5hVV64/c32LEGEVrd8lui35iOdvfyaOeklCJeDEFfZ/mn1rhjuqK8e62znSLZhZN
GusTNua57poQ7wOUKQ2lt7jB1hTzvj1nX2l/4mrfeNvyhyHT6SWgcIeG61qHA08N4NDPtnBhFwth
vrdKa0YZBPm0K3U8xZhw6b383+NuhPDe+7aP9nq0X3AMOPEnEN30uN4rRrn6CjZZY14zuqCy8WT7
PA+zhxpkt77/qKRju46vFv4uFxcey9QUvXhoAT0YraJyb6OGpJutYI124lYsQXyeh/AefnoFkW1Q
nungLIWMh4PXfpJip0ttQrzG6FZQSFz2PPXHrz1p2+n9GL4tddmo6qfx/H3K8bDp1cRzg9HOpagQ
KIafLSDA1i+ZXhpNamqh4ommy7k3N4B8/TVVnkuQIjJHVjgz/ENH7vHta2+Es2N3nwRt5X1n9FY8
qMsCjUTIkx4BoZHV3A1ckXSKWOE7Bfh7Q0jlXwaZ/X2Uwmkimgbrm9Csko7OilXhMSBV+tXUbe4c
RjDwXAp4LBKPLI3CsWydKB6BT3FN9ugW41Igh0JzFweZwUO++IqETTkKS/QKlv3G+ehqO2wAV+kA
WF6FS31NUtJ0+pupKOrQl/mO8A3PC9ffOmuHi5XS6leAPQm7KjortvBQz5SYUemf0fzKy3yvzXtA
reGcGSZ8BeU6fn+4Eu/VrP8t8Xhm9C6JYiATL3U4hOp4uqv4Jkw2OokL8KM6kXoiZjF40hteZTD5
WQWHgUrAe685SjdKBHas5HrpVJjlE19LVZctyfNT0HyuswHhjKrVfdlPdmQPT11kBYDNXi6BCRgl
0ohSjb6dNJkZKKAprBioPJ2YTA17s+LMheIR2vS3h6Sp8rLQudg83+CkJYgvYcsf16H7l8xg6uVp
Ep8kVkpFNAbWFdj3+qVKhbBaMF9EqUutnzWwMJc5/RW+UbQ9yyfW1eOhBZQRwdo1SFQySKs1OsHO
IYeaVLd6Mjmg1ojoG9mokxzf9o0bE+ioR7ZbNEr+24ATwIwg4AkbM2LuLLlM+oq+Za1e5BT4OhaR
71NGFvO++WH2K9mkFQAX4VLXdQJzIRkzPIExP+QUTwL+yrA38bU5y/LIggMCy+2ZVuDSmR8CMhaV
pcSM+0feDR/1tzjG2GZpLgVXulJmQF5eZ/NKRMAH79V/Zwg7YzKQnHqfibJX6vuB0VNXYu5wqrOd
qQR16vcrQkXez0g8Rye3rtcEcbTwSkfN42LNkMeQ7Xbjduxpf8fVmQUQG3DFo0erF2sn7jcYilNu
twXJf7qsYC0Q7PNHm/Fpa2nGRilvvteWTzLSac8J8nVMHMh1jvf7Npp0xFNsTMxh6OOS/6zRPJuP
qwT6CgT18qK+AGWS6mOxRKohlWgzxyWFbRATuvvNe1Rxrsb/KjbztfwrSLSoFWkR7yONWj26WQv6
e9XLvP3cWTu6Cn54BUgFIHCN5M4R2ZQs0FrsKptSnc79CrvUmqnxIazFpxvIZ3OVSV22xoGBA4P8
Bz2SkiDnsYF2p3JTKmXET2aKrqTNLPMj58JGVIxXhpWCV8u6pP0a1d2WyaW2pG7kVQXeHxZlM8m5
NsTL4+weD2TElXbV26YYo2ubInW3+aCD2DUeQqCUS0myzKtCbEz7XvpIHu5IBhIyWHUXgawOUqks
uBWvg/cwA8UUZya4wAts7WkTAJfVLfG66vbAlw4Yt7SrLJrZCpg4ZhBCuQ6cPSwkpb2i6CkKM9OL
02SVroyuw15sUSzuUiNsqeeEPMhmoq1TY8QPfjmCsKpZQcR30r6wixqc+l8SiVbpK6ytZp58ip78
fLxRkDvOM1iG+UNzcBeneX7c9eOJsMtPrh3j2tzcj/v6vG6t7EY0n1wfiikTrAp7WqXrlFzuAb7U
ZAsUw8ADpu+5L+OMe2Z6vDe+YvLYodwSYtmmfQqLyq/ofiWJ35f8hEaGlzaptz2mjLl/uT91N8Gf
Jwzfv114AipvzFDx5QrbptBCOGUx+2tWt5iVS6DX1CwSZRfsptrkhpACdfJpwqHM/ypq1YoCPvZC
8uw8a0wcGzJYkCgX5UsXu4Y3vhicGN38yAJp7IUJCadUQWv62GICFlGpPwLps8shgfjEPkwtcURJ
r/b+8WdXeMsWaddyOxK8vvSG+Qju6P+g6zntLKXfRLKIoOzKFLm2JmzSygK4/1bPZjWukvajIGeF
XjDHJxB1htatgmxvKfepr2Kh2ImEnOpDldlkMG7h/Os+U2C+FtTs3Zob0gTrQ/A8YoZY+qAUD40g
M9T5IgyvGjLJHxUElNGrG79ctFoxAtwn1eygS8bdQ1F4fWPGXRHaHSdZeMTlW3+Rg8F900rnuCN5
Rdb0dTQeBSL8AsuBvdeeN0mfAcrt5T6THEmLjwkFcMbQArqukQi+wVzQKt1dWzwvYdF7aRVBZ1N4
OliqXsWIj261eJjCRrmn9zHH99yYL+oLwsrr3RAieiuJFTjKAW3ZMQ49Hh2tmWgTBk3/TvYqDzd0
eQRZx6e+I4vMtiExOJWAKgaFCLyiR3QiAqTfiDgkVVKkVaDso3R6HGwZvvY3640r7xZlfKXqCuXH
Bd/icmdAuI6Epp7Sh/EQG5pYzg/k6WPIYCmGyw8jGjM8CVbLPP7vMRpupk2Qbs9M8lu0lusQm7So
xtmW22CYbi22qe1Mdd/qSjSduuBj5AQHnnOm2lBi9NVT1zXavk4bmF0MLWljbHg5CJNGsa3mSfmN
avANhr+oruoQ911JiyUeAKDPlfLaZhScBylJI7m0qLFnoN3rp4gHQC+FYPRkz+H188COhrVdoWvB
tin/tlFNB/ccHVEpkuCRhzFt8CoyafOmweopb38h6WphaX0rZM+N5eVj276VQgXqN0KV0einrirp
wmR7FALT0xnxGPVFvcVrL28lldvQaZlfnK9gt6qDNjdk/TuNq0gI/rj7u1Zhz9yv6b331ccNZ8U3
pZgt0FLCVhP/75drDB86BkcN78O+zOUpBXoc6EMvshW9w4T8KQLFKd0I2m8V/5c9yddtFr9A+JIz
HbH53+U/Q+0ATApIrcySNXNgdcj7hBeBPJaUMth9BI0eBp7Da8a6qZVIiy5/PC1rovYFmPRU0L3+
kt6kwgtoEYvnb847pzBt1no77YYCcZsHNUUDKH1HTUICMAoLpmgERUbU0MMtuWEsp4+G5VoeWvyS
J7JH9luC5ENi4iboEdBpa92tBjsvxRFA430X9FMxEdB8RGOQ9YaYph+D4dwf++MZYZPGJ5U31dlk
ElI67i+O3sfQmNP88cHxp3g7qIPLFMsgJZa6FtW3g4u9dDYQEQxaOJnwyTDesnbNBXVmthSmcGTV
/ue7XSFFY8kNBiVG+k/T7FmjxlSVqoMoIsYcmCrn+Pxij6nlTxMaHwagMldG8ZOY7IPm357do4pH
GjkvEjs3c3itjZnyPYEsSoD50a9C/y/2+W0btPaoLp7yjYdWh3I4dsbOpIC6F4Df5tSBpxCCeOGp
MsgXXtODZt6hFT6GM/jxhsP0I3VhwfmEQZdhsbbhzIiHU/idt3i1yv5it0aQSkQYz11If7PcIEn9
AAWudm4NpbShlcy004G6aSOWWy59cGRAidqaaykmye8NPp4Fs0JuG4isTF8LGkH4cc7/Pwa1uwRj
nLtXGSv67t8zr7sHcwyikx3u3kG6AhW3fO0LMnhh1MHB/PoTeJZ8K/hgRm9pmsRa0qZyuRyjRe2g
k7r0blzNU30Fh049pgqvrJJqgdGXPuVM9PBXqZK3L3JhgoSD/HmwnZcifvSqWyMJUgdha/hPL2lM
MDup1cDDXjy+z8e6QBbg+Ovy8c/9YBAw+YpCqp/rK2+Z9gyjXa/NSp1UvTR9V1H02kNgiRqIarQK
aRMpsB9YUJ4Haq9mH/pA409IIu00XbwlMwtn05DYFN8MDC/rimH93vDZcTpSjpsp3vXOavmrh+Kj
OLZSR6BHJQJrM6SMH+Dm2jFIYtgs5Ne0kSuui4AYAAMial+qQ9IKT5p+mSY9WeektoUgodL+40IL
LiN4PzZt0hgFg87AyYXlNXyxjXoSPyX4sntf87gduS89DMgz9vAZ3LD1fE+ydaRDEtRW6YQ4Doc4
2GUWqe+riKmmxrwsO8tWbyhPuOBt36PTpsS1Fk/n4JBWlm+ltowoYdpB8nkkbyoVvjKY+oVimnki
J66tGcbx81mcLosQAJkHuZzdKmPCv/N5wMtdHNKv0KDD9sYOALkGkpWmIrGmXTAJ5yVuIJrwUHlC
L5/2JTXWP+pEtsUx4laAYJBG771S/a8YPM6/Bhl27YnlspR8gY8jpc0C7PABZlfdSsCPJatmL/mX
sycq257ZanrkgjLL9ZHmzaUnyk8GyxaDBA3NiBL1IxEZpH/e63A+poxRuiLIfLha5f9s/sE7CQK+
zRK4f8sla+KEqSff9A0N0e9apymU8INqL1iZTqu7Vj/b9rwJ1tgw8FzkKGZzsNHzqC3rVaEEaHY/
XChmHXG5kZnhoWHu1RMKdp9fq4qid11e8C4CotcwREsrN7I13eS8v6pkqcYsplvY7fnZL2JBX4eH
FoAyOYVla8sPJfpducjkNXzbT9YHXEqvFL97FWTYFZKdkqSELL0fR1RHHddJ+b6O8t+h+cEjR0qu
TqML17fIol8ZO+OsgykKOJWo/g/+ZQZ7THVYCmNfd7Ni1jw2N2ibafZC0c4nFNpKlwASctrgr7wQ
pY80C+otehdph0c2Jm8H1gVf7qzhLaSe4ra6y2sVKbumLouueoZG5kNYimPIF3kY7HuuBxIdSStq
g7W8+x7kMSOpUC0FhpsHNxx76Fog3sgqqVRAzlgRh4th8C6tWYBWPePWTbhlTujgWATNEF0qpCei
1oVg6Tzb+rvnyQsNQBXiuBB3SKjBlQkackBBNs03TQj2+mu1T76+WUuLYpCyRy4xkacaG7CxONm1
j/lBDr3vZCOFEfIIrarNl3hgRkmmbX9qhUGx1PiQL8aY0rUpRCVVjyYL4qiF2WJo3rOtp3yav04f
p459X+mV6OkWpFbfBrxhlDaSLSVQrx3tLKCZx9HN6J45B88lUIyr1AXQ/bwLdM9y25SJbJCq8RU6
zUNkyILiW48WOOraXDxHfd1XqJE+hJM6Kx/JvxVZNduJP4yxjYZ7Owht+qY33fbVhaNfu+zvfgtv
fM1rwklvIH5yOuLIlMoVO1EShwZx8GvTlJLpCn9bKYy5FLu7Q+y6TpT0Mefl0aXMSmqzYhrCM6gY
N97A7E8fDEg1VJuJC+CzdF8eO5XV4ycrm8ujVBqZgR9rRMAlnu/dRyqcK/us3YMKc0DMR1aA1wkP
03LH3EXvsCmioqSY7E+yKkJNPYdR3jHHMVqGnv2X4YA3pMJEje5hBv4zCQUCPK60l1VAqqgLtWHR
1x4lz5/5sJcknlLfrG7ZQ8CGCpkxyRVctPzeEt0iOK3wmrUbW0avBuZCv3UPi5jlwI+TcZJNeyF/
hB55K4idZFo3kTUI3PSKVn4FY+wdStSxXELgePZOjE3rvNVVZkB4onscXH+jSi1VqaGj2NtLqjWJ
AL6h5zZltvXbpUA0nJdFD7P5orpAf35LYNAjqICMCz8JYuslA+0mXM9oX/feWrOKwYRqV0z5OKwX
/qiiRnZ0W8QJPwxLlLzlBIL1vHWdbyQTIhP/v6yS7FaZDM3+gvcppmfiTozhB+b/xJ8H3iJG3R4w
Vbw6LW+uwecveD2DDJbrWfba3acIX76Y21C4iGB2d7N+htWbUq07/J7KFUAba7NvpFJ3ESFmdLdg
F0UUDwB8KBqCCzna+Pb1GdscyAr0PjojXHIb9lZ4rsiZT1PYhZDfjfi+xSARpZMYld4k1G7QVhMW
O3PuOop+OJRoGNvsgs5AWoPlF+0gvQuxKkLhozrD/rCc3X9SDlNI7gmD77y8cOVXqXX6HJGu3Kbb
9/bzV1eUCSsMBkHtmu02DTJKBlkUwA40oNEQmgUcX9xBmM+oYelzES/4AbX8IB6nXOB/wWh9gOuB
+mQYpD9+pAbcNLDc4CzXAcHfKZIUIjSfddQuVKUEVOInauONbAzht0MwOT4qOr5ofyZu5WO2H0Vf
M4t9O6pgQKC4JHvIhP4JqwTylK5XwDhxVFiSw6BfpwF8T2Ttx7oeeKqtxC0O7YewuXQooH4SQMyd
6fOMXZazW+MzaVFtv1UDV6xNmeDFSjx1rqG22TDeEVjTdu1jAyuSnlITwtS3gP0VBzBKboJZwOLE
r9pDV+V2efVpRbD4g31nKzHgR1ppIQABygKyaHnzj40NA9gHmEfCPcI1VoeILaZ5UzlhS6e8NFYm
diYqarKFG4LamS4eth7Zgk16xKkcmOcvLH+19e+tNCjXjCu1RYkWvFEvZryopLo9yTb+mudvQasp
bQ5y9FW4tt5LHz0s+dOSJBjJ/9xdH7I26rSPJ4/RZhUXbODDi5fyStfX69/jV0tC5S7qAUQkyfik
6czWkej0ZOeknoNjdRV7zshS1P9Kb5CBawFToICn9I72cEtDxs/ySeCRW9nkbQ89sXXQVX9ihegu
J2Qhk8Cekiy2t2bxNQSDrbcE73OjtuxLkOQ/FtX09Z072q8I6+RvvMrs0kUYO1MRlCv7PpGL0Znb
ySUfMJIJqsTbcrdiN1wCpM9PdjQwzHFNoZfvBbxow2ISh63GDBwprOdJrXxOdwDDkO6hmg3sTMG3
a+zbqBGRh8y3o2o9qEIKi3t6TU0h+syibOW+iaU4wl/1LYrb8ZCx30aSzSQr4CbmaWcxYE/XQOeM
dNzU1m/TmHSBTf8q56PXqJBmeF6B+4gZtRQav/5ejROjZpu75qvUwncWoupJHL3XXavQzScu6DWb
IXvsMnClS6DdfXQzzgKjx4Gd1PZeEVv695We9hmqeyFs/Ha7Tj3U8d9McvwixLKq7xP+IWwF9Lze
fEYxCNs50Yn5oRM262VwJCS2wWwfhg7V3PtVW6LoW6uInkSpRSHtbQ1XJSwALu7DMaVfgxrHm3cL
LfUHmwHzgtJ271giit5RphIiSGg3tFSCxLvow8aZLLSksqjgISvcpvbwCYklzKqa69ZwoenyeKqw
T9OgV2c5BDVUPrgh/zufVCiz4Yuz01GwJyzE45wvR/QnaEy227rdavFtULd0wpZOOzW8Bqs/lRsl
99Cs/aw2/PDTaG/rwncrGO8p8hMJihBRqL1ywQcfcG4b0+vRW2hBDU13mywgR6K5H1SqsOkkK50N
l12ggMJ2mXVL7pKBQtOrYQADQlwHi0jcRXIUIMWsBWMXJfVUH6xtaeNqxTEvHZTwWM6CZgaT+QX/
nLJwJmlbx5ZimkdShIQ+MhX7gK0agA5abqOEa9blfRSuamrKCD/kxSfR93JS5aYxgwS8VFcv98R4
6HFtHWrjwg04DfSyylLJRNTIW7DYQFx8y1hbJ0z/t0Uuf8lYQTGnJPE/u+yKPUs+obxbq0chTOoC
sYSp0kMVlP+Nws+hfsFFGhw6jASVSd65IzvE0khYdZcrJcm3TxTktGf5n0UpsWzfi2LBBABl/I+4
sKdASJDNwWMkt2KqKI15c1MlGzqmLdS/tBzRbmiAW7UKt19JaH9GkkEqT9ixHtWIlYtll5v/noUw
XubphzQA7f2NIpe0bLyN5G5efxVaA+RFxzRE+42kxxPGWhi9w9vuWGJSttlAy93KaqzPTCS1CE86
TQY2LJumTDFABMAboyZSiz78/BXJTEGl/+elx+oqrf/ExLqBcaO4PCwu62HkzFEumwHT8ExRgwap
WLYdV96kEnL44HGt5LUMbKrPsGaFth17drA68QW0zoA1J9t43adwXsX5jroRASsLvkgjR30NtE/U
zg3h28r8uVNX26EUcxfl+dUgR3irQn6x2UCoZY6fyKanKmO1YhMSFU0d8vLyn/X+vHWMHZ2z+5HZ
rZv4TmGRSM3x+dSjzmsygBfN6oof7yP8Es4FP+tEmhmlEcD4Y1HB15Inrtb6LIpAyaLM3dW7PdAd
9Wt7hZMjbxsoojkonKSPFjOppiX33lUJEV6Rk1gLFVNmVtZSu1CES/y+r2R+eY7QHuvD4GERJwam
FuKz5LIjJsFSDusNOdy5R1IV2rXErlDByfFQmeaDIYhJFxrAu6TZxm00WvrQb75us+ltgLvvGAUJ
bjEqXNZ0U8ZRgQR2pCjuAIete7cAK2sfr/oEhhDL2OST/4ZVjtBQgVjU7uB4NUgbaylAm1W2UBqk
0MkfpB9UovsVnNmEYZPT+YmYFAxjTie/RiBOUPuzkObWdIkk5hkKu59CvOBcOuVqX+6qG4eYPgNE
wCPp4AIAszGhuJknodbOzebzAYvbvbImCiQrOAxqUIeiUis5PUPEzeBychml6eVx2nyaKA1eqUbd
LhP7aT+v+EQ21Wg6UCWzkTz5yG2sIAkT3WYwOwl0oBzekpOfWWrHahwT5ZKDmVek1wwAXSmDf7r2
wuOqWu+pdb3YBORZKDadRN5tdII7mdkOFmK//Ni8VameiXItF110sIxUuKp41msLhZgDNx4V0R/k
QQNHDHH/drGZzxfEp27ZPmzhd+UwcTVswR49EPqecYAr6janNPfuZTX1KqosH4x7nSxIN0LewXWF
cDX2ItgDkip4CGnp1SrTo3BdDx0f43r0vS9UZdKIMiupQOr+tJ4QxoyywJulNxpHXK2N+rTWniI6
8xPygmdcxq1DI3fP2XOzfgi5zB1WG1BbKJGe4wdunuZAvNC6gpVhsdJi0BHuYLlWk/ia9xU0bdN+
8lyD/FI4Eg18CW3ujQbrjSHdHz2RzK/TbLR5h7CgLYr8gc/OtjwO+yYMcs27FoB0UjyrRad/DGbk
/Cng6q0t76XTu4arVxQesTCHvSECpWfrP/m0u2YVgb4nIg9AMSfK58nqMLBUmeb13IKopc9NTfac
JBGyvHQMIxb1X18WHGdsummfHnDpCmfZdFoG6ofe0/hH3HQIWtJWO+aT8fnfbsZfdBpsTwv+MiWv
ul2k78Z6wuw3dzqVyhwD3amKHoBC3gX3u83he+8oTso7lHkeWUeSIUIVPbr5LRgVO9RCCW3GVwod
xM+0xQaxcMAJvc7+pygIrWAkq2t3JXcja+P0kwSsEBlu9IIKdd04xdjX0fJFR6zvaKI1z9OFz41y
svisfp/9nm16mxgAztPCDIqPnGG9lzXjTfV8HxnHFFmZelrl8ZNd2s/f16Sz2nEnSx/u0NecFuzS
0NIfxQL9bi7AcS12+z+iFamFpgMSmjs/Z/Ke/d8S+EqMdeRTBruR4SM1fSW1gYmhnJMsMdR4KseZ
LZDXPbvc5gYVwD3EqNBLyXojw7TyUBxmwj1EMFQpvnvbTwmBHk20ReIgjLmZvAlHXLkl1ql7Ruh2
WILBCYnJ+Gcz/zaVabDXEHQzUipk24VxUj231eJiiYhZ6Cn80vxfs24z3/C2g1CG+iC7aUI1uJRA
rgN2HfleqSwX0tau0X2qM3fN0VmKx8gkianLku0UDC+NbVDZcwT3oJX4aJuK0ASf8nIGiQsXYgWQ
fy9D0RqrXJRiYkWqUYYkfnSxK/59NLtOY4iFOmEQum7MElXvkQd/jwSOLgNbd3tKXMiaOE4a8xnh
KXaCDNiIw39Iq1dAZxy5RUprFQYiW/PZgQzqDmrWdoLVst68L8t40O5eyQOv7daalfPpczH/m86Z
DO9OWrPCalmVuIPki5bP1wIP7d6f0Y6WI/wZ21mG3aLkAFPF3ZLZngBHBw88NS9paBjylDUUZ32E
Vcrvm7fEHfkyo/Z7+V4kjkN581W/D+2oBhrrax0NX2iJ+MlrHdc9gXFHtFYPDcYRNLyKnTrptWfu
9zlhKf14mmi7eg0MgqJepAZAMFRbtRE/qYq0Jx1G3PZ9dDnjGhBFcsfFaOu43eNiGKYDOM+TOTtk
wJSfEIbtVqVfuogczTbr8/Udjmz/qJZVtddFAt5IgKXYR9OLY2QOGG4pSArrCZlNxOFCcyjVbFSg
1S4WLB8twMEomSEUlyD2OMoj6mYINTs/akhBwc0Ahmc3ZNtFoHqSnldyx4zBAqT+VTU/mEArWF6S
iQD69vHs4x8acrDk2GPvxTwhvEeGfe6HVi/iwKPY4NafQwPi2dXuOq2aFWjsd3/HIry+uOH6QiKG
T+qMvztFNy8bnxUc4A2AEi0Eu75l61yPD2ODBab1a57ItOMvFJxu7YkfrbXOxAfrxRHxzFtMSBOC
u9fTthjHvEntxO+rhmDRMQgnm9hAwp4BzTOjHgJAlY9Gyr7QIjXwBA0AhUslPLhoArVfS0ucP4oI
0L/l4mpFiM/evnFJ82/Lx64qoM2hnpcM7b8QsMjh6NGq/xTfNZUbL7JTae7qSbZ9uN5zDkhlW8Fj
bj+Bs88nqpD2El/DfVUg1PF14OA+m7m3iJftDHiwMPjdNou5i7aF9Jlc40NlpQ4XjoNjCFXwtl+c
XxQ6edHM9N5tXP+CY9g7VJI1wn5bdhJOaqI8vXd7eoTqvXTQ3RpJZ1fTuNrHm/eCBbTnwH68hHLK
Mdu2Mpqc+pb2cN9r+XAZ4d5U7qInhePga510GlfMHtYKOM51Rp7uV50Qq+Y6TSFEWth2XBXvQfVj
IaWbywaNDeEZS+aiQZAMCaE+av9l9++oqXbpdavUww36k8fwxykjLGHIVb1dTitiYgrXE4KCVknR
wjziJJ7lug6D16bHFcCxiTxW/yM9sFZ+X+vxQpNR8Tz1jplPgFXQtp51t9Rf19IHPzG4nrdk1jWi
IwsRqvQ912H7hecLUQXd/3CulfdvFsM9Spycsz2lNBixKiS9g04ZkC5TNPxXU9WicFy6EWb6u8hd
QtttLVlMbyJ+SK5sqDqD5AKMjrdWOOna/oaSNgxRv1yOVZeyjqWwMn6vLprgWKXNlw6R3mTBlf0v
ulYwZ0lc5Cy1rCMiAdQ9I2xDxwcx6PMPirq/EgsxYuqxuOMkcvwg1uln4WKEYOPUrgPYnEjxapzC
0bqZUcFpYSV2wQGrVetZHtv3dPT9JpCV7xlMirZh33LTP/IxajXsDF1nmFpch5BGKEfvmUuG9Sxd
WD4CYsnzBER0VVThBAlnIzNdSLkIn12MtzcqO/WaiSxaXtl4+uXyFamU/vmbkZKV4gje5gcl9sYH
ePd5IR5lbrNtMWQzmhM0k7o1PCqhgHZU00z678jfynd1hvK4XtrtPe6mNPuZsN0lUTmiJR9flkf0
BAQ7csNZoZ7d8w8Pzdk+RmgOESHMiK8x8F9h015taC6D8dPEcb8iCg68zDwCTMaysDffZJzKX+bh
II0cj9U2+klNksKuPhYRilgAtxC1tzJjJ0L91o3M3Biy5FO8l6vj8GeWSwR0fRoUdszebZ6ygPX0
q3LIqYJJm79lasZMmk2daxCFklBHHD02kQiJgC8lgnckccwZXfvlfumlOeC53FkkaClzRpFfn4au
MCVjDhUJEcO4d66QhL2qolAUqBZTBopdDYFe9jLgmEhBKTKRw0ZEwyTDf8pIlEr7BFBKpMToyjeK
oifJeLhaqnGkYZ5h1A3fQZDwARbA/xgyVXTBWD7oGu2eRN7zLsrYqMUPI6wMpLgsWuPmY26j9wHE
FYOe6RprWdgiPLEbx4Ml6AF0p6CD3V1NP4FEBl/Wr2zVe9IBx0Etq7dxL19uV3L4exiU59lz+8Qi
/rqWpMpZqW8ndxl1hfRdT4yICXiEFopBMMsPyDCKfdHu4avye9SJU2x7ozPTd9wXDjFk770jp43z
Ik1Y1/znIe4h8v//psV4TjdTSoV47rbRp3i6h7RCcdxPTn9vLoGg7el8AM8ehf1gaXbtHlDsDHIn
ZPjXYUARhrj7tGF9Ivbv7BgSaISIkTVKVgmY1E5l9ya5frJTB9+swS70/6s5SazY3bE+5Rpye/0O
aEsyLFbPOWhFwj0wRzAR0GwEzJkI8tSXqsonIA2EZPrdCD8KCKYotLZUdE28MudV1dapLjY8VhN5
nCD6HItuJPdbBLgt0eA8laLxHm9EoOfcMK6LPZgxr4spDsaWNghgOWrEy47qnHGKGpq8DhhNf2Oi
EoDZS77tl6f9H8JLmoqfSHjvuMCIphJov6d9YyxVvRT+zq14kwHu7+M1VV8pWmXX9n2oG1XvzUlq
FlUPGplRBFNEcLyhrcVgN/LP41tEauOStBsD8khx/2alPTjuV66XlJsboLVwR4BcK0ddodV8lf5o
iHNltzc096FglGolkqbULUg5mcnwmOEQO1Yy0TLbFP98gNCW/UhyRL17JrOUmVfJ2mtJ5qRx2k8R
tLjmFiJk5ZnPAqDNRo1KqZKMLIYAE/LDjf4wYs6Hxk8CicdI79ojLSZIQy9CgTGU4dJonmTV2tm7
Fi78l2dhrprt9tCyAmbir1EiFpSuZpDEfYUpYclwLR+O8+IK0+MSg7Y2QaSXVH8yEwadjPRODFuj
uz5/L4Zk8IsgnhRS+Kq0rJcLO7qpa9GVbz3ppAJZrCLrwuwPvDgKzHOe9AMAKubpdrSxSaeorF/3
sONB9Q0rDPCzwrDi1FMG943rMTfTVDQyZMHkKqo9d3gQzuzgvxMcO3J/teP3b6qYWPBaFUNJ4dni
ERl+ulrOf0GR9P0CqxzG6b3EIESZAEmdwloSkUC7Lot7dzE1v90FxxvwDIS3f/2YbVjjEnAuqgvL
6FJ5EfIqGjMJUP/yjT0Jvz3V8dvPZ0AFFB5TEwtmQKTFtsieAkrsSTqQo2CLcbCek7AkVx5PPe7m
PjJeckH8qfNyL2rUIAKSbvT9Ms41B3+YgptD53CwwtWON0vUgWELAE6MiXShmU0LcTDfY4G7kk1K
tINBfHvYWmAG6jNqbsKRqdfSrrUirg7mVP+bOyfbaIwvZzaTeNLWV4q7lvvjadMgwqY301PaVdvF
v6WdAjxIO1HutjKz0zD/fGAlNVHP2czGOpipNc1uji3zCWCTp3+9PHf+myFOxf0iMKhVg5SHydz/
X2D5gg8WnlntdGELT11398c9aIZp6muYkVX69c8S4S9tYGQ4gazu1YPIrFs2ZvBuq9aohGHN7x60
4pZXTomr3BQBClU9jh14wNB8MeAPM0pVcfZZG9ANrlFX7hLRVA7wo0dlPZMCvhSyrUAuGoBTuy9A
D7vyQ6cMUKyVyqGPBRtzT5qCsSDeXUYrYkapmte+Wvaz8/Eazk7sgmMTZ25fdcR4O5QgGmBHIO4Z
yYKE+8ctjfPt9wucHK/t9KWM1OeIfTR8Z5L4ICNkvtHk204E9oA/+N2ulWYnNGDVPDinVY3+qhOr
DX7fIYDhmMTjCViqLjeIK/HlPMeKbLe4tXUZi9HEdrMB+Za3MFLpTrgE1BP3MC29SEYTNAFyNhQt
yDZolPambM7wbPmCqkutbHw4X9ePhpGpl+D01ozT7Rq+Cl7CE+fq9X1frodxYcfexO9PSsqmnb/x
stbF7u225JoHariADBMpvj2IynYpuKTxFJ0k0GA9FRLWUC5PjZ4pkBd+3aRvzoXgU/73Ium40G4c
qE0X2IJxTVr+TkDHf7vo9ZHbkzzKH7dQDHY4n6etnnSHcol45A9Ek42D7KqMe2gwRSpuGETtDLcI
VGg6mlZfl+tDuc5k6ypu0m9s1Xr7r06IdnVatYZohOmAtbLOrgwdywVPX4JaMADd0kPaql0sw/bD
locSpLI/ZleN4MUstKB+BVRMIga4F9TkKO08D94TWebgq4c+L0QgE0P9uO4UQ+GEtlBCbzJsNoUn
JZJqQWWY2PpCWvDutztqtQ9eKdxwXDP9cDshVFhd4rW5xz3bCcmvtU7gogvsuOzwD1ZCdGptUZXj
QBt7Dw8XgWrHhdgXhax8Y0apEsIJw7tl1QdIfJzq+0HZpnpzRDUiR89usmT3y8YyVlvBirCOXBpS
iAy9WiUR8DsZ6p645xuRf4NDpzRogtC5eN6S724jOHMt00TUWeLc61qWcqsNbZc2sXBo+iCTp2e3
RiDvak0VQV489NWS+Wjn2nTV9ffRqAtuRnoe7rusonblqm3SUaU3/Pj7ts+dmh8xlHgdQIjcHoNb
oDHxozjRHvoRcHfPylOjGH4NB9dyHLeMapmcF8tZ5glFEalHyQRf2tF1C0sr+GRu5XNFLFypUOjU
pDaUiwE87QG7sfGUj1qoTFx2K7sa1+zc/YtqMfqaieFezjL1hCyCHdMTXWjP5D7okcASFemqV0bt
Oss88v9tnmq5CTgjWarZ+sVBazhsXcdCIRiBqFegeVzPbbOwfyT40WUYAcVypNYFEmeUZswb012M
GicRBCMx1KeZlk32KKJ2wQAdM1EroAzpVskgb15bj040hcptn+kKyEEiGTlZQ28mNbYjuIv63l7q
MbwpvJsvYGLd+Z9pQuLALmbxELdMg3geyJvhSKnAr4b46pT0bu2KKo5Wz9zlS4kTYmxiwqQNuiou
RTOkWgdYd/j4H6PkYBcYb7NcpjSB5ozgAnDSh2LX1rkXvdIbqKqwi9k4+8v1/3hNXmnMRk3ZN2nn
xMLh6Z54IzYwJdg6Y7B0gDrSR0SCa9OYAi+5laZXZ+X0b7LzZw7AIbeR797LnxlFyW0gBNjOhQHv
5bocDgm6EdNbo3oiKm+yIhqSJWMHdk6Zm/rNJXm8vBUcxGwsVXL2Wyhd3smk6V8Am2SLumn2ZBmu
LPk1NIN9t/uEt0QRnC8rVQ1zktnX5QqJb2jQGaKjKhknHwiw5HomfY8VxnzMLiwP2xf4yoyR9nqm
FbkcIEKTQvmX60xmffRP/wJdGR3A+ySgOS2uK9GlXv3kiqXOknxL5vYE8NOHtlRw0ICbQmOuIrAM
JoKPPpwUKSU/2KyamrizPlO+d85D6SAhP8Ec8+of/2mQzOuAAYe3K4Gw9kN4ZZklXoCWgU+B6DUt
ROTwbi5hjh48RGtv3k4QWVAFWOcb1G+iTerXZTHEqtMZ/+1NYyLhmYyFR9ufa5jcka8zKCRG0jeL
B1X9STDv1ssjsNtiuPm/c30T2ix4sY9kqb24aOH6A4atm+25fI7NtBT9AFcRlCwhat1LwoS601vh
84eDdqynQzRWT3JHMlXCxy1HZwIMDDEDkmVVQfaFODMyzNCxEivj11i3n0w+YsXBLTXJzdelR4tK
5ssACM8/Wp74Kpjum/Z2gxkDdZddCMXYHeXVMuGgVgL8QoBcPjMZedprGo+nsP2bd3hZCOApf2cn
0VxjMwt9MakoO6FZo2rEvNMMox1og5NsS5076pprPgtt99rr/AmscQtClWhoxnTMIXlyL5lNKKXX
ZsgGMRyZ+wOc++VqSgyRB/wEVWP+y4mbs5XY5F5vn/42rPclJS07sbm+Y25K0VsEBnx7b8xggNwG
ELi8XIp9CvkTDfthVvCuDfDl0Z8u6pWV7E3g8FhH4spFHt3/l4qkXTUCzX8L2yKAT9OfrUbmjRh2
ImsFD9KjCchSd88sNaaLDaKTyyksVcUCHxKy/IzxH9bf+WaNMCPZXbamBI/Qhe2081sT3PQGosb2
Tgea4kckK2t5wSwilOkNM5C8TMq6k+FjbVb/4pP4804KBjHZE1qjcUKiw+z31MI3BWG+vwUkL5lS
bKfcsvnonc4AzHoanHKpQhHRP27z0pu/nr5kXUgCW48WOf34I3gadljxwib1NviT9hPJawi1ryg/
GO55IWjW10CDo48fUOPaJiRhVum9EIgQeoYXFgYSsQMSkz2IRDD2tAiacRiBqGUUXZf7r7aNHigO
x8SNsZQns/8negPjd1JJ3o9VjDBkXzHBYVG3eQ6C3khbjshWvf3CgzqqKF3ngPeRbDoIVWGAXmpU
zBXKxBM/3lEGGx3Rp5DTYo2YM/sq5ujMErJYp2Cy2jUaM7VIXHPKTyNwseYeI5kFbxmB4yijlmvz
mYloeOI9DLGkim9XDTIrrfObY5nvxkpClAUbph8aA1jBdzWyjo4/TvVybaPFy7WMmmeSIC1Xkox+
pcGL1JF2m9X4pa3JYE2M8SlUqJdXOC8WSXezhKa6rpYNozaTivTSCGM0j4jZfd5nkvLsJVSjj7S4
g88RWDGb5yyMXSKpIkyfXWmw615RiTC2I6Mma+lsdzBo9t0ante1LYWpPNWnvZRDbxX7B3+ou0xo
4hN6R6jO7KS3rpj6Dp/8eq6eSgSHJleX60VnoacB0KXFN1bnc7Ek397IEfbrn4tnT9sXYXO7FNmg
q7jdvTkyky/dNAMRk1M3ZQobeAnkX1yhSYhn01xiqahxOM0dYLaz9FMUgZde+bIkNRtXiWSDMTfP
BtU77KZUO/WSVSR7w0gm6TJvHS8qX3bdcSu8rnYkivdV3oeRfWH5lHOBwm/SSZTVhpLDmrPjYyGv
nmqZln/4hzrg2bOC5RXvxG5Fw1K6q2OPr8++/0wRcvcs1WGA0Dxb7SUp7TBokgEuhZLR60lPt5St
NIvbSLcrG2HHW6mwvrZfUkZOiZilvag0cdWiDwM2G7SKhBfDwLxrLkWEZys/laZatw6fYZNrzsiF
2iCTj4up5l/DiOjDl+sPkUQSvT/RUgXhtyPdfN3PoV57kjq3mAdK38Fy7pyyb8HRLp8PqLd55/4H
bHCi+RAJHtTWFuChYpsce059GE3k7ZcSHcStD+tnG5OAeFUiUkNyZPp7FetdzyTC7SnTo6Eu/zA7
1XimMEwOBCBUzyDW9fPCAtiXxR5KGcMrcps+3br1dClbDWBS9damVBYv48LQZPTEIMFJbChgBVRj
vtC0HCXAsAO5xm/gNBrSnX6iEgL1DmwpX/c3HP6nArMrZTym06KuH5GJw2WOKvVaSzMzfLSZOHeR
7LRbXytf3+gSiYj9KLjPAQpWc2Y7Sq0dBHhmGeH0R5+jvmGjzquBn02ldszonzRnWEDt2cBLTG9G
LzcuAPTSJOg3mG2c6Fxq2HycXQBRLY305o410CNv5AAsnQyl/+hZM4H83cBOCTo3o6/nzvSsjrhH
Nk9o5UkClKhA4nt1ANxNUzrHelh/CDprqtfKp/ge240pgpp+Y23N8/7/rfJGIkNUuq0YXg3MhUDW
qNIjwm+a6rcHMxUV+EmYIVlMuJssNq0RlWMvRCX2Ug4b1Wba30iSWSfYO3YVxDSH2qK9wlAe9mkU
lHH4W2PZvoGvSH9ShGpynODfAakPEo0NtoxKukzgd+EvPTp5096kskRv2yCwPvg5EXJ7j6fuzVGQ
u9vsRSnWivA/I2NujefoD4AKFI04yx5J1P3iF1RWx0PtGG4HjQG1ZuYsqdWEY8D3WEvbnyvoNgvV
pybsl3agAT/L5INC+IrTLtDMIZDQMnpR1RfxRxHyJBsdW6qgxb+mtR/muGnP43ELbqZ8TVOFqcVE
ZBI2Pr19rCAgehiDqoev2d+YekosP6X+B4I3QCak3BZg0JFlEOS1ut2bNVuHv+MQm6isnK3CG9PM
LeBOs//759Q9mY4FJI2H7MfwYEaXKcZW7h1uAZiHFvq86sRsrkuO7iJE+wpwEggiY5PEJHdp9+kp
IS/aKrZCxuOOyUWcsBYpL4GNxz5S/5BuXaBYz7w6ToHfZbuLnCr0tl7JgXGJOLFMcB0xtZW8o7gW
DI1nVogYQtiJhIIswKwoyNljdBN3BWRMdZvdHSaLW27Likyg0iwnwTKNOcgPLBXkABddSIGLWGq+
2WVQ7oYyfdwl3lXEVvZSVRFiNABa75Ocv0fBG2yxZXD3D/h6am/ffoQOYgCDiCXzrw8f78izquAP
Ry5e/8rL18cPtnqkMqMdid6GSyoI3PzfFivFfOCHzFcvBydQgmeXiq8+eNTF0Hb8h8mjE0TZcZZA
HosHTT9h+qcD7uRzNFJ/qnEINQGHGFuf+NjFkUuEtwk/GkMdU1rUMbLqrJoL2OaYDJqLqc/qjLAX
WZBxG60b9lzWxwB3x0uuMiDDLK/vDAKsaAjOWk3OvuJVx9bo0H74XQ0u4eJLLLMuoFcP/iHp3UTZ
Ha2idymP9SdFOmOKh+p45tqXSk3JKVeRioaeAz3XQMiUUHDgzKVyNOBBrvhmirHTD77MosSKZMbr
W6e9cgSnjybvnRwUrOV2fw0iyZlVeYvqmESsIwF4RUP4cZFX+biI807ActuuEHgI67ozMbVgx4p2
Fyy+i2Ggx0aOZrqxZYWfYY8mMC8AMlxhau9C73Nkeuk0FDmnj/eOhz1IpiYWjmptD7mAivH8Fkzi
cFqIDZuxl4n0E4qtwxAN1vDFDo7YeR/poJQKfkjdBM/hPXa8ydNKB0RX8gxrhfz6VEnmynWvvKTy
3qITZBCllfztNfpsTEXVjMLamHwHMKEoryL3Yuc/C/8jVvlagl/92y01sMdMzgj/3KPCcCh8kvri
EeOdWS6+mtdW1vzn9Rxscpx1ujJ1KSIZS8MSmEo+g4GJ9dd/iuNqIhujeZSw4OsGQEYRzUZ/v/Ri
FW9sLeELsAqXezjlyAgan8uUyDrbdHxzeYMEfkmuYxJZRSi3AxgrA3E/J/r+WfEjgnyNw0KOAp1v
fHflU07Ge1/Xe0qG6+WJhwYscCGc/dkqfvll8QqKohCps1Xy8TJJatvCXcHhP7pvhzEwew2alNxY
iszon83X+zhi1DLrI44AB4EpreCACezsE2zysJCHPUmkaNm63Bm1YXFSe/xmTEhzORRdrWzvKovB
83jYpmrnzdCimvdNa9QJNu38quFPNJKOhcZffapfE320RGI1qNWDRj+Mni9Y3ukj8LYz+NxpBuOl
gzDfb3CBz+H/EfFGUIftSbADu3BvEMJ9ypyFUDUL96fh8vuCcNkKHf3gJrrT7Kry62RBw9vuGqCI
zReY9F0m8qxe516Fv5iLm/BW9EGgtpWFq1tcJNoBa5WDvwxRfUGKxxIRE5+vN/DxSnweF9zXmhZU
Aec4ewuQczysYtDnaia8Yf2fUWlkHmF/ZWGbhYg94vj+egUXnKwl9VPec9YDgM8KxljOFMQCR4wB
f31km3088k6mLhdEjchBOjdEKhjBPbgpPn6gjMS7f6bFa7oVgQdVz5r86QgPhZA6n/A4bDxTalcV
gR8THazwzY0Q0xw6m2zrE3UT/Xc7M2mtjA0SBGSEAYeTODF9AQo6lwJ3dq+n1rH5xB1uwvqFPqS2
Y6Jxq+6XAqeuVlk/jarqq7eHjdxC5i5Lm0yp9okWa/WcSWA8EE3LR6dnRZ7TkFW8JjCyY3j0Of0Q
nssmAezZDG+ErrSeFfjfy0Y3DDLZrVcrK1LDI2Tck6/2fe3GHJDYeYLAaDKiuvEg9xmOeG6DkPT/
XQLdivlAGbxCGmEBOSt+5SCVbNGSQ10EDVDIi8h7T5EaXVi5TDQwKU+JK2Ktzv5JK4C4IBQ8lHGU
qLc94Yr6H2tDimE7Rz0BE5ckFvcoDQTaVTzVNavOUCPOZbVIXeeZ63BV8x0n7SUeJ7Qo/ksrgUw5
2ItNU6bcArb4J418ToXs0yxQe5/NMpZs+gFbx0XHDbaBVUqxQIc0eYkEEUZwrz9Ap0ava1zrbTTS
anhDGv5V6ShzTVX9oy4eZgK7OK+KI7UIlkPvJcIAMeRLmDZkgCNC+n7vCEXHTDuM9RVtO7xsZRW3
ms4NQ5abnv9VodA5MQys9LrS7tpEU/qnSaCEHRThYPH51wYw07AOmB5LfRqcWKJVgmjAtCLjyFpY
MLLEtw/RCeltgypWXkm457Mj4sPNs1DBwCKixU5TbPdKPuoceo2P/RWy4mJTbjSWUlwKdAY/mek3
pN7i/JeOwsXSCLsUxfTt+BdZmK84XbtAjxtezx8v3ubvMCG5NO0irHIOFbBCLN6Tg9ZNO7Djo0Es
wt+yRqKLZG13tpGUxW3pUPHGdlWHYvaTFW1wvmIth9SmlvTw+FWbXoCBhk7jhPvoSYJgZi1mEcfj
yEIXUDz+4ZoDQl2EERKDQQNNglI1+V09RuavNQjMl4E7DmOFB6PfN83oEPgq51gqY3khur5dNbKw
oWzx9dHpgzz1lIfMAKFx+ZlgkS/OBpS7LrzsmrB+uP70aKPI9h8b0NNZtiKh0avRVVjOjWHzBbqQ
k/jewAmonzDNdRfNbWnKTfXClMl0MrWpcccmwpYa5sk5wjcZMQECiHR9j6I9hJSDPvvG/gsC5thh
QPy1BIWrmBfBwKKQy/5GCm8u4e4baBqxp5PvebOtT4mtFcCQav6+bnBG0poHyluZDN+Y0Iosa3pe
1wImLCpuaAy4OKcgxDF9oS8VhSOeoHMjPv1Lba7FOPz2tTnvB2VvjrGSTkdN5JjmG0PbwtavWJQ6
Lw5qAP1UFrGo4O76PYAezsAFInIu2fa8K1n4C4xTwqUgz7Lj0N7veUpD/XMParIqJvXyhz6Gem4m
/e2ARw7YuKVzZ1L+Zo4FK9HrMqE/nj5bDS63YHvQBRAmth3/ATlI8HZ/RcdGPfrDcl34Mk1gyiLZ
RaULaMbsmTY7EhRVK30s0xpOkFyiA9+W0bKIWmy39nZp/1Yxws2TeSBgzzNU4jsuF4SeMSJhP4Mf
3UYQxQJO9runw9UJPIBDZ1pBztQJAxNSSLjyB8B3kvTZbh3t3Dy+rU5fsNzOfKJFoEIK1o05vlUf
j1ZhkUzW5NLoLxfNIVK7GuKOkwlCn+6lA5biV2nzDlV01wNHsoXo77xKhT9Lt0xd1huQVLudABll
2os36KGpo1N3P5LFfDqyo85dtZf38mNQIM3FOuT8VNbg0QPThtgF97TuZ0EQKpBktkywj2O+3niY
XT53ELQAjNV/fWBHEZzhnnFZRRqFzwfcySKBILpG82tN4hZgHcVAFnVDuFf+r1HPjnhdAcOJzuUg
d5GulS6DO3fcsEay1rDk1FLYu72ysBmd7KnzUUw8K9Xve6Na4awVkaGKPLsTpmnOZr2hcXFi4kLv
QV5Z2fjKfsn6LHR8ZJtSEcVvC5i4wFA64ECu1dHAgc0yfJ4ww5ZGj1Np7ICSh9eVkmG0XUp4+Qh2
yTzElksf4piVDmdPqcqRmhylImZKFN2PO5wb/+NdFabkW4SGnpCETFxR7WZ7J9dpSahCu8jqo0Qz
gs326kji98oPjrt8em/Ot1JOn629hoPTJMOM2JplX3XPTSh2z7G+5Jtfn9VqCe7dEXnqFxj6XyZN
Twsyh+D5dQEmgiEtlrvUAD7FmwITd6fz9ypXf9NwH7nkPKqOTPI6mwjjX7bXeoWBAOSjR3xXQgqt
iknNmVZ6n6Q0b8N4V9ET4mHpJBR2CVskBAWPu88zimSWa3vswCxFEtKdFpa2MFl5CzGAitwCiOSs
yNo0lhx8iiO4pz1nLypJhfw51uo1bOMFWPmpDOGfzMhIDbyruw8aibHvhC09AgCi4PyuRoqZrFn2
S0U6v72ywzpmiaqpwk3iQ/VO/+hYdUC92mg8CZNjEKXS7uL16HdM6/MwY4ld9rrSOtCu0lZFR7Tm
KoSqGfHGK/xo5yi+/OyX/778eds1d4H32o5Tfg3LD9jv5DkhhtObmzd4LXsrJQkgPZ0NPXLHhXZD
aKCR95Bn+PfB6FGn6+ywEcqoJbutDfw3FPddjhufUfrfXYrbFqJN3oPPodKvhYzGXLSc1Cq/TUkT
/G/nWPWXCgVBWpdMhlF7NRuErqpzHlTFZhHZjCoLUHLNwkv43cSbhHgQDiM1GL5Wg4QVvLyAkvVL
IS8JdR0XHLkaLMc+22u/GF48tVJglfwPmYrsFnNdDQuuExTPLmYm+gOmsu5+eYfOLPEh9ysNR2y0
7LPOa3iNPviqRh4pM2h1Qdhkou4Gks8pUd2Lkf7qYsw6p4LL8ve4pj9UVQf26ofcnuuYsLSxMl4u
gJTjEV/x/9/DDCG1aE28kiyJXwR13K9KsQt00CXhJKr3d4XcrTCFwJ9aqULVxEoNPU2oN1rHnK1c
We/IZcz9AsLeGMKT9RgCITFHhkN5WZWC8VAcjM4wMLwjZ18cIDReqc19gewVsw0f1RQu1K+OwBWY
G5X0dvzwC7L3rmRv8jjwkTl7Ng5SzWZ0h8zB1ns5AZtTcCHhaBmqgLosSBgcK6hRMvTXZWJw5XTJ
90/S3/mbeoYHS+Cz7AounsJPcxsNYMjQ9VOHkWVNxeEmasjQCOTQ1Ik/EKUgN95r09N2iCI4bQS4
VWJl2pOFMNu4XNhprdZnj9QLd+WLpzqgpWvorzOtWOXmCEW579mxH6AcZ2T/KnP3EM/WiawpZ27/
vCCnUultr1mXRh9eIc8yHz5tKVAtFtVkCXIQRsVISj0d2UP7mgKSf+go2FNFRD6el63ermE2Ahni
s03tLV2IS4Vuseacii4wEd+4Wk5Fywp3xabm7FPSwjACWmcWp0msdjDWfdgtDnVICMB14KoSJrRm
JWTVCv3x/GCNa/788lHH3+0WpqKk5o+mjkctLvTH9aPO6lbjXuKaL8bHpAB/vkBPnq388gvwE3n/
zPIg3JX/0uNEft4I8cIkjp46NUuoTD5hABbS0q+6onRHJiuN7PSw8sLyysRZ7miVYYao0FY3J+3p
+eo4bFF/VV9h+4yk1OCQXI3QBW60tP+0b+r8ojfrzwXAp0Gub9w3uI79S8D3rRXwA2JgT/A1IOxg
l9irgawsGpvDOp0R1x0QWVx0ocWdclX4PbrM9ACpF0ILvtxqq5cYdQBHOomb2z8PePCCSMS9cJB/
7BHe6SU/F0Q24X5ylm2/ZfUTrVv/qLIRs6yOrpLZxIDGyAfyVSNOZH6W6tt4FD3MfmMHe3pvw1ap
/IPjnOilCpCqLG0XP6EOS6en53U3Mcv2sbOZRwReLQlTEK1Crz6AtCx87s/jNlSLBbLuj8lRsw4O
mDaZF7UEhVnO4yMeLZlKLsDoIClwneuh8zLTNV/NO9jXe2A6gmhffEHcXzNgbRrhZM1s2FGPWR8w
jGa0xv/3zN0HdgjPx5QPfAGLItuyJkoT1XxKwTDp6VuhMh1b7VD/IMTw1GdZaM1ZMJWuKufPKC5n
QI7UNWNezQXZhctpBYFKsSBk5c7+/sqC/C4HmTA0RxwSw+L56GhW31BmXb2zPBe8TqbuAIoCE2Xs
CigJ96ktpgHIv7tPw7tQlnlie6suaNMiJzbFMaoDagqNVwXqQV647+iuOVL6atvU5ZSu1Uv19czN
hMrgPYAB7BTWq/ci1/1Te9/eaom+TcYrxSRiZ7pNlo1jEaDy3q4hY5FRGY97+QQyEZjwQwxNejkd
JcZA2LF3tAYkjaA3fZSmIX8pALKHOr8dueFCwNimLYGfqPOl6EkK58OwmhOGoVS5PAMzmAMiIOD2
nAekPx8QDPwTUc0rvQg7m+aJyj1CUeD+l1yg5D4yE02uTBsuRhOLvcy91k0fDdRLhAUdETJkNwmj
srTNQgVdN2fHQkdkV3bLA3skULjIxwZF2ionjrT7gx6pMr74MRhFpk7D4lFFzIcVRpGgLAeMeUFj
H4VgwXF3jygcNPgwDxCg/midkdxS8AhsjfSamOc+bnd50sW5HdwkcNKvwwNsQ/FGJSaHjShSlHW5
WjlwIFuO5vAg9YVYWq1GtUfT0P6YgwYJvkLijc4pOwquFIb/NNzjCuJuChjH+zeHDl/U6Na7kZ+p
X781Ydd96QVIJS1NhYa+e467hGAIEnAmLvmqc6lC4WOCLiRALEqRD1MtlqA7hL5iiOKQQzdAgvIO
h24geNLELNANxgn5Hh7Ay5j6EomzINCUPuJrcoVI/tl4qShS+50BCm6WgtulOhCzSDTXlgyGlGpp
W/O5j88dm8BHa6zM2is+/ER47AVCBulm9H2MT65sNImGnZlvLe30KuCl6Bnhdeiz35oOebFxYwoN
emurahy1ZLH7HoGJqzsq4X9MNCqJAiWg9TKn+F4sh1Vm54zJ7NtUCUWE/uXsqksWkkWzY+8k5FH1
HQAQiFrG841hZKWhtJkEsQn8l7RN2N3xcbktmN2ogeFgJJq2+n+SfT2b9AqJNpCdr0F+yXiIC+PQ
LtP+AeiaD0cZCMrO3NVLNMRdXKb4UpvGntK+XQaqP41k8XDp8/omk1wagDu5uathI8Qart4H5I/z
Pp7C3NXegYLG3sqOf49p2aPXfLhzvbGj3eN2oTwPHe2yNl2nm17puvzPF8MKx0kWOZfsb1lwHfED
8x8dMpivMJktEo/n2MGOfulCrF1PVw/8dB1ICL1mcIFgomrIGrMfdnnX+q7n8lEU9kb5RMb6GmJF
10fSqTruG2fSGqqhjyj7sJV06McunIvJ3Yze0l1g6EzQzA3t9X13TSXCQMsEggoaNGXeAHh2TDti
AXwdUBCUAwzSAa8uf8x0HC5fqMMvqOrr/MExSoRtBe0fAhcrCRvXqhuIdCAZchkyc4CxWXfvaKtr
KseDAr7FrHvVYSRPSH9ws7uFBpEuJfzbb13hQKOP86barzqP22g082J7wI37KCSeoHLIsSUwJvcC
RtgI/4xEGoFSNMS45JCnhq45nzdwQ63uNbdkMdTJmApGfsJilwcoQasrf4gNSgRUMjsMdNXMuLtj
TJv354/li+a6vhphEbxkvNIhyg8f5ueD1ahdWmwDxDdT9qBymVuo7VrZOGd3unU9/Hc24tJ9FNs8
nRgakCIGO8jhSuV7aVXW6o0Cdb2kYJvdtU8Ufcokjh9gDYFaEyAWreD2+qQvlomtlzBKT53g4pSK
sB491MAlKH8OuUWEczleUunYeAE5oH77BWV3DwM20MeT1oKv7NI7zDNlvM2xdDhu0v/+4ctcZeRF
4dLvvtsF7ghW3x6ZCzGYkscESwd8sWH6s4oFuW5adxzdB+qSPdfF1v2+RaPpiFOwZiRAP0LJS3ur
nY4xAWg+f5r1RuBeu00tMT482LYRly8G0E9DxuO+eHHAVBpsZ5R+FG18VKDrLwSSlq3FapNkOlSl
dpJ5JHBp5JTsEeSDBdl4GhNaYRY8tdKKyjprvU8kSYzQ0KPMnXlbgBkPEhBJAz0P8Ejc1mMoXTit
5c6IYTZmV5s6dcyf6P7w5HnttBRaPREj+OnvMqZV6zesGJzV/LQQZnOPGMld/BKhtyQmmiPtiWXw
O44SVUqN4n+oNUC4V+/nkPEjMfMQHkAxZ7o5iiBYdx52n/dtHRnFse47ai79n+Vg+RQfVe2Fz0IR
YyvIx2iYQU1NzV4dEYZ8wbM6mLKZacbjGG8H52u5IMq5g5+fJuRop9UkCNAZSSXJmswu88hnhidz
DOnXmoILJJJQMRREbC2lT/gmgeswyKrsT9BYrbDUtPM4zRfiDYed6hN6vecn2Tlm+QoH5uoydLVm
PPa4Ski+JiDUwIH4VvqspL2gN3BoaQ0clUKNFadmny67yp3y2CrnF/4ToviIb9NuDH6b3Y3GaCLh
wBoMuoSan4WychqN1E/Vg36c9UAimQDMnOaN5ohWc/dLNqSkjCvk8//6yx0qF9GjIoUir/GvJy6j
auD5gYGFdnhwQEnkwI7a0j6zH2bUnTqoF6Alak89clf3aspF7fExyictW+71pNcI9U6mqrD7nVrS
KZQGnu8zN/IicU7V4Gfiz30WQ0NyqqF+u6nCx/46IDGrn/NR0UKi8or1otSxpKZohyCMF8SdotZS
Y7vREdJTGl4ckhxqJ0m1o8PLeVhGww22JRyPcaEUowIT2CnUnEIAh8NzPOai1cKyOu4nsRcI96wo
KboSFckhTFwU0A1I46+HiZ3wez+h8AaP1wwGZWEc0h/eGTc5R/0RPYNNDcYdCIiYXqO2/rnrZ9Fl
OLSkFDgqzaWAYooT/sK+AzpBpGpVlBsNJqeuaczP0OofJ7Sb1HdEUSpJBPanTKyNO3w4j6E9W9WD
F7HoKWG/zsuWc7Ox7aEkOOmSM/E9Pk3sbsjjv6iYEC9+tnwJhWx7H5fN/+j80lfrpHiyWmXEiXsy
PTruH0q8/CtaC0eo1PdzZVjb7Quf0N+nPeyAIsUw6Br9uom0JtpNKiOec0hpHkNInTQiGdgZWGTv
Z9M950L/S7rhyYNJsl92q0Xfnpf7YxOoP4NO1c3E4V9KumfW5vNGdHToPwRknTkKEPCNEsgLHpRE
iRkd6hDE2StUw/mmC/zm4SpwhRccX0pp1HKxQAjnWqRq916lOIWkzKFE3+gY4koBT98hEtBjdhuS
igH0/hAfvYLlVzCnoFK1955qNkSXlLE7jCx2haev6YTJPI2xltkMR8dcKmQ8aKb0HI0J38QDN5Rd
MqJjr++fgI7ZA8uJ/WcGd1QqEVeETSw3HHx8CogQMNC3s9zEAuTM3VIOPH/QZmBWXjT65J8RsuQv
l/blICBrACjNiuYOUnnP0el4lEy6eRDcoGKGo/qlvvsM+BK8cqWCjl9spIsHvcr7RpEhKHY7qEPQ
OY1xxGaffT4YGd81POSBuRKCh1Vt53EW4INyyJfFsPIDIbFV+lfTHjPErYKRSqVq9mgzijfxkhYo
5PqRqjOTuyEd3qXFaZcezqE6hk55vJLrr5e+LwcXlky4hPIK40TH7+jE8TwEKMCHBYUBaW52PuYV
+viX2FYXvQdZMY+hgOdRUQDD0lWVorRHRL2BPZihzKHyBB0yDrhV7ATv4JLR78XWzOHlCf3bww1g
+6NquDI+YGO6yapiV0vmYMECQXJJQfX8JZQYXRkGByLMDAwHBJFYb9nNkk0cAnTciT1S1uX90Ozo
ku6evcHV+uoAlZYbhjj9pf3ANEs9RHnffqbcyQVO6Wqj4SCQA+Fokfh9++jFUtK+B6L2IAhD3LkZ
yc36KhsNOXYmyRsdTBlVsKKy815z9OP+Onl3+/Qi+4PbuLm/2S5G1IA3o8BUTqAdcAXmclo1fxtN
dPWarSx1z5ohultcLKmJq23SpIcW1O/LvKCr2iucwKs+ICCZIsF3pI+crNL71vNYYeIWGlB+tkx9
P+Dzg+WHMkbg/7NZzSdZNKyl86QHnqqBy5NsI0vuNOIvJty1X+IKvIYitRkknJzkBNuhNRDHIZrX
qq3pr//dMCqm8ymHrbuO2MTUHJ/wDZJrJBSLjueanDn+C3AuHgp9OdjYko3+uIlkj5IrfUZ7RW5D
bKxM+D6Z0r6cflcsDIiGbeG/BTyBbnTHJstmiZB9NnDVHslwh2Z+I+awTpqAO2rdW7OCHpLCULcb
WPbQVjifjN9QbOSGLQX8yjkzlvcYO9OyOLrV2e0GXCfCdaliF2yzHe9pxqK0aZV/GDjp3dY9c3qP
w+AUN/HaUidg5sFHBKRqPASWH/l8HBFst8SFvK6WC3VQVqLj+/lAIh4Oh0CdRm1rkbZ5Hq2y7HyZ
i6HXEMhUI0xRZj4/MyN4yzBLNvaiT6O3M7SwUIbku9w74Gaw2pZHSEWxMi8FYS4vR4cs3T2aTxqq
mn/lc+97Ioar8D3iMmFNNP7MhSq3py96pQgyUx9SeHHj1qtEY+HNCOk36SXUIpHU7NXypltd9q42
YbhX74J7dr2OJmYERDpyWVbx1pBbTqBnUVDUsRNBxFgrtrSwYxWxCcsXecQfYf9gL3224Mz1F3ZF
gUvwLSyYjrvqLKuVrPu1D+UAJ0Q/pm6VsmAdlP8M4PTI/jzQZ3s0kE7kjdXDc4JIsuLBW6QXw1wn
WNi94lY0PHg5Ij5FEK6YrvBwSLU4EfTi1Um2QDlOCR7xBVRGehYPJ2PWO52tSmqNIWxaVAwOOjap
CSBKmb3IPNWPAZRfwnEBH5qEMjbn9q1/z/znDgAFHYS8Vg7FPaun5uRstSEn0r7WDC8brzqDCAOE
Nl2isqp3HUG2bTkTCX/L0PLt845y3YUAX7v/oS/NyXRxWbPWIWSkkPpzvLOQxVHMMIS5IM1Rrs13
husM7nmN4ZYJ0Hs+2S5zKLgPKrCs+uSP1hPhvao8BEAWjaZI9beVvA29DwHiia5aC3ZyVZke1186
HmDZUsg2rISrnbM4G6yKUDDJ6lNj2Y8Hgopbjl8DNFX4gq8t4EEtYzWeWJ5Mms+IsD4VkuIfzIro
XaJpIYryLABumKhXFCxOcZbQyCN9z/9VzVv5gMyq14quyy8u5yzPAxK/7rfdfAKBu5eMGeOHmITe
bVfYuHw/BLNqKwt6IaLDy/EOHZgaQZnSYHkZ+EKzjCdeh0A/43dbkb09HzD90qB8O+vcghfXdStz
j9xAXCFdfrk2qKQzHTjY/DJnLS1iNueJY34OQiPmtDTAeEIDgZOVKKfE5gAgdzDhbg999YtPQDQc
FtbS/Slwnc1vo0pw1UtLCMTq/lwdMF4hh4fdrpKLVemfaFWxyVnoA31wMGDB5u123Bi8JpUdpRYi
TVGGkRJnyriQSGffCp+WTnAE6HCLgB9scQ/XFZ/1TrKr5m89Sp4ZFxOji+O8n8k/JG8dhjwKf5H/
4ffEmHQTeXen+wciDkEHGMT411D1RlqFLHuAebm89FCrqCis41r7Z3H7i+gSc73BvF/QVeAOb/NX
FN+m/5dKrRi3RIc6k9Ef+ena1O+G6VG6BUrhc4wkBPSk7Y2EbzvgDx65Kvwhj3PRERGBHvSKbPm8
YDP0QaWYBZAEuyRAPHLONDzOuqz5E/yIVoHGWf4H0EzBeLjbvigsj6QiNtl1wSDpCq3u1snnY3Ii
+LCeFqN3KRaMYYJ/3vG7in8c8rjT0NJtxhik+aaR8GtQHlU5kg3g8xE19VnroKqhBUBSRo8a2YCx
X9e7fgnvl/D/I5N2AHc+zVg+z+L8kkNmYDoo34juWki049uOxfGnvfb8FLS82S26lx2hBRyhvcSA
mkeRVBO50wKMkqrhWBfu6CcjeGe+Kj2uR+PSStcwtg2miY+CX1R/my3aD27DN27zpQ/aoKP20KvX
tohJYyD+zhEtkXAtlsEYj4Sqo9hMQcvj9TSgU9itBrk9W/VnWFtBiAbPXl76sMsNnXoe958hDlYO
OA7/dm8XR1fvqJzoIulLrPOM8p/a1szTproSIMGYeA2SZ23x0ocGjnzRwrdpLPHb+sT04/mWlfoV
jbn5tpV39G8Q7a+oRgsOIL+sJHtbxjilI0nyhFESjtZ+0IhG7pM4esfPwpYrS+Xdf/aYMW18CGLq
sUgfIYBiEql8J/iFzGKra1ZcKujJs6CfliZrZkCPv2iHN3P3dZupJLMi+pli4zNBycb4S+h+l8wS
filZBbbHFkspex+Jkcrc2fpRZ6d0oWGKN2hwXW2zR5FVkJayI0ZcvZYBUA9QozyKhq/V/WuCqf8Y
7j/1YsHfdmxI8nBugcgawUgBAwruyEipMLimsWg+3+mcLUSM1r2cK4lh78ra2Ftenmrs1X0WnUph
K1oDQVP+MHf34s1IP26H+MReoVjp5iJunQrnnKpZFV6S+msISd5iM97JbkXsalKibplzzv644IaO
N497N5wT2IiIImzuVgOsd0BjAAdGxAY4xvnTkmt0f2/mARUcHEIKJZfW3UoH87pxLozwvD7+XILT
qBcBu+Sdp9XIH22qVVKPM/i7+NFhKar60qglVsBB325B0cxN7GcfQ9wiLJCkHGIWt8+JNxcAAvOV
OJLPhMd24Qt+AV7cN+niImCAhLd253pHmCKAiRT62CalL13UoudC63nLsJLwtPlacpWzThyW49tW
57QX7V7myR1VGRSMrL2Twhtk8WHkIAc717vJb6nAvIZnEZkiltEpR+t+4ci9Pm7ofu3EonSUm6ns
1pS6cSPkCL8HauO5b25xl+OmhtFtOj6wXhpY0uhH02SKAIroUqIlwIG1NrZcysibNnpeKuoJhKcU
Mk+xC/wTns0jCANZ0BBRezGWp4qfYC20e3DG1HzqVZfvmyDoa3FloWOIpcv+WFNGpg1jjJV8uxUS
v/BaNcsrl+aH7vyKo8rOAG8Uw3FVZnpJl1tsGSvWZYttxi3E0hYE79sddccjZjUh0BdQ2y+2Se65
ebG7MjTBsNM1NPqtExbeIynwhBvLsRj5a3y6633U+Goq/beeG9SKAD/3avl8WWeUKji4YI3VHFJl
BaCTwfXCtmMdRYHzyRez5oJcX7PMZGIEiofyzvg8G0I9jrTFBIUIqHKIdJSIl0RwwxymwckCtVM4
8XE4ABKVxfjFpMKuhU568l+VGSM2/5WR1ZTgCsK7CsG8yNTqzJcAm1sjeaPCqQkbnEQraTm9vn+4
p275Uw+IEVJgEp0shGLnVjUQhIx8WqRUkx1rlFueIHKfiUiVmaYJv17a631T2rJndPgJ8QEkoYu0
1xrKLd+6iY27MF5FpIHd5KW9h83lHOTXaPnyavHTLZTjosma62RmfGDqQq47u5Fidl7/bjqDVZr+
ofnBwpT6x9caH4n562NOpLshF8v0wuei8z152grI8wOJ5185pf7WiI518ObqxrrKMnkLJmjGJZ85
Gzbp3fBwU1enyow2luGfGk8ZxvZasMZVdlLn6Uf7ajuqdwcNpbYNX6UEAMPJf/KB54kxrx4UGu4c
Egi5n2v34h1nMHm2smWLTxwJSYtsDz9+cnWsebWP9Fmt+WYlymLJqY9tQ1NgShDwijwmsl9c8PQC
tyyLXUs787Ni6swyw4BzC9XzX4HThrdAfSefR8bQkHUVzXcLuamO2xx1utQcHUCvNQe0GXKHyK0O
DOwGyYuMyyifKIvDmYEIYAg/pfMUMwvD1ttLbEccfeWiK60MxdTqbwKplFlc4Y5kExgCpzcGJ67W
Qa5+AapTRUt0wjjhQSFtCQG6baAVoDmTKHniPBBRYDGE22BscGzK8bYvF/QDgO225SE3EIt6LbhE
VPo2MXXC2WB+aMvqLOf7pF2Zy5Ps1IQpiTen8MIWbNd28ukHUc/c+oeCDR6Q+IG8e5c5+ggBklbi
3AN3EVH6Ha9swqIugSLalUW7QonqBkvX70BemqIM4PITE/W31l/xKEqiaNQv4MT4D3mtT0RpkcEh
85LP6KDEMcno4M5Gbd2LfmlKtpnSm9vB1ZTqorZekWKrb0kWgTRc/pZcSJB7AxA1kcwHdVpL5oQz
6AqEJ32xFTUf8CnLsm2hzDXXbI6DHP+fJUn4IUuwzn5NxEk9mGmPr42TDcBxjMlqxfa+Z7CXMSrV
yCYi8p8dMJJ7Df299YxBD/Ja2AG+UUKFOs4kqxTFyp84QHcGtHiUPArLI8PyeUCBN7BikR/dm/ft
ZG3JlFnnsCNMyATZ4j0QECtDG7Jto8AtPnFTRVbJsx7NVu4NE1aOSK4jRegMZ+jxrjnRrs4JfKfq
JvWY7ymu1Pgp2vNKpikPXInOpnizYXWzfDGKCzvzCzNuhzN/fWiz38uJ6oqBS3ktGw55j3b/P0U5
s/YADAevsCDLhYINnsfaxDsLMzYaTeYUToNp3bStKyJ6B2QQCwrPH4hMnXSdoojFtGFlGfq4A37W
oCIUJzqz3y0nttIsyek7HaBdtvVPPOfbKA9cWhg+IGK+aj60zqNbSka1AXjHgh9xNDGzs6Pk1Wbv
xx4pKFYcCKt7DwSNsHzvp3JyV5Ju8Vl/Mdk6FKa/oXW7Xxvq2tVbUhglfASOlBdI+rajZ+gK55Qw
06Q9LEXVZx0B4VLA7gGzPfqY4cQZnTIuQ8hiDrYPEr0cyjyHZvxSrDs48E5tvwMVtGVoa5acWEc5
IAAM2f5r4cQJSrl4q3Y8te2XxShMpAjqHgmyILn9C2+6UhZ+x1M1AjDmq6uRUieL2xtLb9XVJrWa
MS1ojIJYknjhoi96HWA5OBCfOwUmSLYyvWHG6ctZJbO/qOcTV8lEdgyA/K3veA0CD+H8/SASYKKx
PwZmexgxx0U5BjFARvuRTn0uuWdSo1DLa/BEZDAHyQ1MnYlEODa9KJPWF4LXBbOgI/pbSNge7x5O
3cokhtKxD+piAJ6DlljLNz9MMq/YOonfxjgDM7oxQZ1R4UTMk0lgDptOEb9AugKflnjzVYvWzkoZ
ib02Z+9NK/5uP59Fl9JyUrZeIaw5d0bP1NAZI+G8S1rEQ6LmYJ5IIThajYhY7qMtWXOv5ICFFvgS
RYaQYYYodLzFHbQTvQCZ3BenPHArdqz9Ww1CSCZjf/IA+OZvPohdUF1Zye3ts48mz+80IazTR7Zl
h/3XKZOneRuqCenzIMLopfIy1wOA2FnN1Ve1pgu/bVtSWepgTQ1JIa7Dlh2u0LXDlpctEtOLUNaW
5TbMPsXFINcKDPTc4B96GYNsLL/mY99w6njeO7+UMv+1dJ2jau9pOcqH/xXeup4oBV8BDmvzY1Bm
NA66QZVlfEIqUH4MaGUETXzRMaj05t3Mm+uRjJtTDYbNOvZ4kxd4Q+T9Yz/KMgZK7l8HTrf75jxU
bjVzBH4NWUIwao0YtI+C5vp1s4QT+6RuXu0BLKHTQpWYfxk4yLkEQCOo7GR+WSe0nirRibEmWegY
a/6emHSJSh+oSl3EtaGux8UimPnqGedQjQ8bjoDwY8T+Sn7Dd1GbLkTL9gRJIviHrwklvM7Fn2CL
+1Dbdsjpxpqv4D5QvL7LNAkLRc/0LPEkhEXd4VBK59VxVkAiKgzbtqWDWQCY0mV5+0n4PaCxrqI5
oqNKCRcgDAeEd95EKFo4VZbHAAI9w6tApXu3sIDafvXsQ3cZE0JzF/P1Rf6ZGTY2XK4UqU9YzSc+
T9rcaApfQcaD0+IV5no0XK0ea1k68OTCZmjliJ8hml8sxfCu6L/c3lqigTsgIJFylOoH6zUb7QRD
o5h3iU7ApmedkUmvfz5xw5VtMRORdEvhTpf+zs9jb1N41GD0HD52j3uz99+ei71pHjDUpcvUqiFE
fvOC/MT5LXOZTU3UsEBEtAVeSqpulCtOVDg4vKfBCp++mrSj6N/xZCM0ffRGraql7Ppl2abnNoVu
PfrAj8zp73z/jrpZVwjK7VC3znQhn79KPgXEobnaPNNYUx4g2eNa37Eb//H7Pz76fhF7+noFhy0t
het7CVQyWCcmvGKVRvJ1SZbNr9x2ZFwsRl/8PKueyp/laJvCeWR9se5JDkowDgB6jKbrvHBbwZmG
lCkT3walPbVAzEIxMMmXSKaVfxX0GQCCzrMzouzVfH4YpKLbFuDV3yBLNmZjgGF9avfFSe8Pho/d
0Tlr/kG9/PdiOXpx2lDCcwxzvKC1HQxWMR4ULTWVyoeYMHZDRegmbeTlaPQrfVp4YatrU+BJzcGc
HOwNGUxkmvAeTMqCY7qwsVrJX4rY3qeypHp8dUc+aRCVLNMtkVVpnIOKR2EoBUxagHG23E0fr8cG
VzFT7MX2jp7diQPaC4PObAcA10E5qd/bbVDlSKekmXXndaAO+6JYR3XZuh2Pris9vlFmKL+KhtSt
Xa9BkBr04JPKadKEOWc3bsuL53sN8xrpoYX7bRRjgBvuSUCnMQzXjKghmbwxAMdhe9Z5WaY2TnEU
twecFfKMPgjKDpYakG79kZl+W0/aA+byhqE5bgssf0uekgmHGQ5ArKQbWUUlKGlDace8EfUlfPbm
H9D650RkJ6NiXzNoz9J7ouqXHY+fYzrWSupytdyNRDrWonKjvjf+4jIPIUb4hAvOjJszw3m6leR0
4z+VF9SkVO/nQX4BDaKv9Xnv6GIw7HP1oqAvoko3yxaOuqcvu8YdbH2khdohsM8nCLtcr4vy0KE5
FcVWYzEvYMvy2mZg23Ms8SwzPG7bswKRnthszCo6k7Iuy/qP0zh+L+EjLlLiY7g8fF0nCbfL+EEs
Rug3uhCtCxNk0qaugZFrYV0BKyygtR59GM+RIXYrc1g2kTyfoptb+scljH85k5bz2q+uDoD2VcwZ
SCfUXc4p6ZQl3X+FQsDuDfpWyV71TZRhtcYBaPU5xlk5XFOYaqAPF+TR3hUMhzW26P82o8JHD0jZ
xy+OxEMiam4Fq2goiUQBvgAWOmOZqU4FogxXmrJ0Meqo7AuHEPvsAcIvc+SFXK5oXpIBI8h/OVAj
5D97J5ozxRPW6u810wPpwTPf/NxQVxmpatMfjCrzoGSL+HyjGjBdqgKJGYJPDFg6v50oir6I4Vwp
U8tWur3oUtBw/5qfpbgiQXhK7NprKjQa5d46yHUWExMX/8dhqthtETYrewvN83FM9Smm21h/R5pg
ScuxKdwjJoCqDGhB60jHDXpbDX3F3oQHppNimqVzBAsAZURCyb2a0lR1zQcgt05g+l7sSBDek/17
ZsMJwuMIRk3thlAH3sQjxSYw9570mfE4akozFJSPXF+WefZ3xHFNwMZDwffkFV7fSisYwZV2iPDG
OBjX96mjmTR8tEoKZbtr99BCix+juVhXzKOP63SE//g6W3SCIchg4r6DCXiWjJGgS+wKc5foiafC
KzyTxB0eRDKSjkfgIDcNLC3xjwR9akp1dtPDGFv3Z2xYy0xtmQG+7aUyWRb2sNdU7gEsBpX6wkHp
mqQbDoHz79tXKdU/kasECSKFoXaPWGiD6uKFWohQfArytt9xv16HCgItnx0WiorZZASsqFvJLBR7
DPcKaSK+xWqrd+sZgMekQYEuM81YmdncuM/v0csq4hbYR+ubnme3gqUHJRchQuW8BK6KIXu7oMYN
WfV60hBH2QRWhd+H2fLQFP1cszijk+BIAEB8tDfrRK2ME9eU3YN44dKTXdOvCQNcTKe0jIq0maHO
+U5a0nnien3HMa67G+THtrBZI4G+ATExgZffB3YVF8anL6pVKzgzhAFYNOYnMmB8TrD6lPwtAoJN
OppiY7xim2tyrSeYKxriynyvA1wLzPuX8/NJXIxxbR+7IiBuQnciZaGuR5+991kpZOl6/pUtp1JC
S2loaBK/yu79TmQA/jMk2LMhBsmqLRtuR0rtfm2SLk5T4DKAbfKRudO8tBsDJTCmZXPv4AKPYdSf
6K83eej47i6vlFx5+H8RjJ7GW7R3eAnuKb0X6IeZ8eBEaLu0wYJvAHTJzfMAoho/uT6B2Jjl/aXe
7TO/FIr1WMdZFsCWB98I7OHj67i632MBPD/Qyi1Szp78WdixsoJAkk0PIptg1KWhxVsNE6xxLJLI
y6XuczXee4lChoV5by8K88+opTfngqyyby29HNF4nfkvXZDvMhXKrHxxORIlWhNs6HEF5siygsGX
iJp6Uif4tPCtR+Lx01U0f9K8NztGmmgBkCavIIwQwUjSQYKdR1/dn7VqKgKmC6X+bbzJ4uP+dak+
pmNjgdig0HjCos1Mf7FGJkT4AyTLPINJLu2gCiIZnRHeFQBx0xsvJsUTYXbpkaAR2J9SnbtdAZxm
WEFAHVGsQdrXyRrr55nZYf60kioOd0Q/apQurNwE6iyoF4h2KsloPAWXWf68mD4qm7BuOmy4DjGf
ZtPXh02TAzBNPAwEVZypYmtQiDtxMBbpKe8rWkPZDLqab/JKrca818jDwPydLQHFxQ/v99XZOwvk
uhQa86hE5YzDf/7N/wkojEB3usTbasBepHAA60rSxyznSlGt4nEN1dpghVxQe2gRq/zJZ9lhizKm
aYDV6Rzcl2o7vlOVZNAZ5bT/7r/lqmO5NuD3Y0cvJzlIsgu+ONlIErP0VzfoCqg4Gd7v608njnaG
Og6Nvf7yculmhs1k1bEdY/5SLrB/gfkSvNUakGk5TIQ0r4VNhCy4Uz/MOXuRQ20cznPPZN0CBg80
WOudnWIJJ+h1YDZK+fzmsrLVfut4mHdOnBzZ+1LxqUJlppZMsUmsO0ls+fKozXF++QKZ5HXZQxaK
rnXYN5MDSvLKX61ir0zxvL4CcmR/KE4WioLqBIUHC1qzgLlFYrVy4gjppKQE8QwrX+1/bxQayzYC
N9C3av8mw/eYrubdQXm3O76L9AVyHVDCKXEoAiAptM4kX+wMCUeo35YmHMRylenIScmMZJmw2NJx
nF5IMMZy+Fj8EUQJSpVh9hc9Dms5yOC2I6Gmm8QPJjItKVScL7GU3kKQ16zrQf03luqXndUSQiAN
JHozXuBkEzJ1XFDvLVXclUsEclNHcYY1+C7du6pBdTMuQngSBFN7/MVq7jy+mkbH4utb3iDwfzZA
+WULpMipeVY1bmnY4brnRaTZXBkgl/g6dMTzswBrT7MlWMcQ7S7VfTa119ty0FCHi+kZf43lK0UW
xUti3AjUoJEkxCfttaW5oZbI7zeti8Jjun8dURyk9q7TjokwuWPxO3efSjE9B8ftfj+vyX+3ayjM
1KOKF4hnporyCT/mMf6hh97j3JJf1x04lKBkRq5NfWvkg0oDhnb0/GUGgzH9d9Pz5kQYl6ciquSA
YhhyXwEsPrCmYCG1pzHt607SugLeZTAFo9kzpoSdBIO0fcuYikd5DjHbgnPJCToMqFNAFyEaPCQs
eafCOapo4yJ/JgCDL6mo/buxJzmRBxaCYUEA6SNNoDXMJ3SspaKrzGtT2UFlgRPQNbJczum0hk/M
kQnssIh6j/5Ug0NnUZi7PWBAQ2Ds2JIZ3Psg7476FSsHZFPuyXY9Ix+NlAoMhE+MR6auyBDxaDRT
KW6dK6mnkfn3zjnafxAiOpkysMyjtRx3pDMq2ZG29yfU6pqpEB8Vlcrrbso12L51ddfWIpeTjCcV
+ACpfELL5x3Q5JhesNnKFhwEqwyOqqCozH7khAMq+iY5A5WicKk0fqjrRU3eUzJu/8K8MqrlckZ+
jIai5yQa3vr3ev13O0ePZn5cfOBq2z2RLgkCYdCiG09GFPKYohfnMcDC/8/K3Y6Gbw2JOC/WGMBZ
mrQwdWCRh7OJzkdXQgqDNkW3LbRFL8e0I+gq0uZj4EpAzeYHHxvA0AAiEYS5QtKG3eAmG3eWJ/NB
le94W/rJXMSHWnmlCBod+9nBQoJeTp6guP210rBJlJk4B483Drbxb2dANGDkamVUEqfhFvsOv9ps
6fPBGKqrIQvcfLzz5nidtS6BFgWZk/+6tij/7wtOseyML2n/u8Cy5fajSEKMEX9pJpTxGCuZDrxN
kDtLTD9ukpXdTyIOLUGf7suzg00t9dWrVtc8da5wknQO2j7/bzngyzeFdWf+4taB+WEG2FgiUkF6
574EK0+A0DMm8Q9ZAYjFDHPRpPcsFf29rfefPsc4jCfnpV0ME7g64AqXcLIH5WCBV27jyymrjHzS
TrH1yMMpRVkFJwrJey36Ot3F9DvwLzgz70UhxuzrQeMqea7vvJ9H0VgL4/O7kMrXdREp3A4TM+IJ
P0ARuCh9G0Zxp+II+XgUQTObn9yU7NprPgGYTds+gcO6OCJ664MDtRKyP8W8EC+VZCueJhPhVPS/
ACThQzd5w/9t8z3wrlFQZEu06sAE6nOnDmCLSKVbzxYLifXf8Ock68Am3EqqoswJo43eh3b6VFg3
lYyYltsRAKzx1pQ0JjPUJCxcnbPaI04cdobQg3cNPD/R7JrRmtV3C3UaAl8N6bIeyorqHQlFTeQw
gyMB9U2Xoq/XtVlViz3ISBryjgyMMpObxVkWtKokDnqq0PrGcNaC5Vr7oaIL6sEMqv5sblY8zcv8
HdOHLWB1frlC7Dua0XlSframGXyyTR0bSM6hkvYsKgtBSclatln1i55k1TL9x0LxQ2ZN98i9ntnl
WU3ZjIdwQT9OtGIdJu5BFqhyOQSZbPf3JU06vlawGhRXX7ml/FLQ+/7SRABWVYrCj1MG7mEHGeoN
UMYdEKV+1mBB1TutlYa+O2/gmKD58D+DE2BvYMTX7+2tKN1Xw+cC9bO9D7aD3eOEzfwiLRqUMoCi
IY88NF07Fubnwo6sQdC6tneih/IEL4RZhzZtUx6WWGo5gysvt+t4osWtjXEeZ+FLfwZIpt91BXNf
wj4+hYo7zW/kNQ6f6bif6JkQpwKMoXYwHu4BhtVLPCZQuDrN2ugnSEAlbi0Rrzi+l6liVyv5nRms
vlBSyafI9/YqRZYnUew5EJu8jAV2rr4hDO9jXF4LXzFnf5rCaNgoKxqdFP+B5z+AZprGdMWd4DNu
dVRi3/zQMz0cNBsOjScisYPW7gAc/8YYy5IHvcsdbR7iOz12IZLJRK4g0vOu5zajOXifI6WRyzcN
tv8tSU5fQ72qb0kMAIfp7I1WEjZD5LQZ5q3dk+LCb/IMw711SRliJ6du+fz4kaS8tI86t+GsOySc
2f+kZQFeFE839cgN8On88oZ8n5ChE29BjeUZHNOHhHQovbHrCVKb8bJzMQqWqmZAvzSA43WYUHJC
egTr1vlo4tja9hiinmqgDLcLkk0JrnIBeuc0U9+AhH7RG68fUpnF/qJeat4l+uhU/f3Rbz1rtXDn
+VJFwuQ8dv3LNDQMQs/b/gX8W2aSrzjm0zlWXAyxE/prXyD/zeRgLKF/4aJuoEFCVskXHHbbJglw
mthCrdaPUhljp6+8dBdPgUXiM2gccktSiCf7uXKOIPl++DcFDq1JJD7q4I2cWZhsqkIDB1IAom07
7vrjaLNXU7zYR5UrbHp/rMyDjt/SpqGsSV0UK3GjIo3iGLN+ZiRL0TUsoDGNtT6tS1axZqPIFcON
g1jp8x6OnP+HkSuJmOStZ81lyOKsE07u5l0ohYAvYZ+FFdm8hOgoSOp1VRN4TBTw57mTFOlGxkMS
N72xZt0r5EODhjzCr5V4tMeygL5VnY1aQr4csRYkPdQNKl4sNwhlbhp7d7ZIf5ogxf964GYu1LA4
GVsb/S1rNzlXESmPHoBgXDljO0RX90z6Olp3ENT8LXqlXDMakElDzXrnGAcbKwf+uQdi+1UvJsv0
iw58pxTiAO71EL99Q2UwQX5ZC2crEExW2vaJMjhKJizbyKTa1urV/dRuQIJ2TX3Aglf5wrXrnhBb
W1TLkx2AqLBTcgL9Ny5pRJsAn2Lu4BQjp55/zpkAvVUVyOEDeHcfar7oKlTGvRro2XxYE11/62Jg
HOQVuYZrZrWLD9ArVN9HkUOLMTqqJ76NpzoqDc65ew1s+P44RrvN92fDjNtvVpUj0Puer3+wKOsw
VgB09vogpMzkNR9q9RiIzCH0Ue5qnjSPhBtRqgE6pJEr3oV13PSrdbZQL1Yh+11MqOM01cNuIkeb
l8BQqzwAAh+MZDh3GQEqGZdh/H2X7G2BIyl9Ngp1g2BjUin61RStCTgZq1tijKKIvTN35bRgp6QY
UsF4DpzomrtIlwJGq5w2XIEIODu3URLIe+Si1gmt3uyulLOpepNxQ70FSrsOC8AEjkpD3WAgntcH
7sHdHW07BWrw87EGHV/CWp/C9vNKg4zWIM2lBs1UHueESCSfcz8SkNGV9kGZnOzx66EGpgcioHug
2JLwui8TMgzHJucxiQJC97wWBPBnBlnSrmmc7lZJNlQv97SDzEF6beSApyBimsHJmC29j2MkJ8rX
OgcYLH5+xKlwe2Y0/l67JgQT/39K9KblDg40lGYkzctXBFvNaJtE93R0Le+nFSpaszUXGOE95ujp
i/XW6hQc7+EpuGrEDf+9LcNaqeUevxNa55oX57hqflhdu9pr8Zy2QMfuxNlKpgNeMHJFk0mGu08r
I3kFz96hCo3Kh3LNOgbFF+BHoZ+42iuUw2yh3SydL6cQDMGF7vGK9zKtSFbOWJ3pYNfbFDgZUxHq
cyvyo4khwbCHWK4Sd/0ayInshr8T9bm/g/bysFA93jpwYMJkJQtdzj19z5VfBFcS8XeBRc+OR07K
lorh6WxLe0gz4HH49k2bxgdrY60FP8xk5cS1T5RDHs672rZ5GJvUS1zqsCEb5tJcOisksB3h4+yQ
TyGb9uXeie5HH+MPFJDVOk5eiIrZYr/5mbtYQWsVjmt9PKLJKgBXDyamATFXrDSyE3kvVnoRICAW
HE+cSDBChxHYoTikXtg6J8MzcACqDiuxO/uoV9LdCCPHNssBUYsoZaXhW4OiBzWOfwfhNyX6uqML
E5AT/xLNT4iJwW+r2uRZf26pk5+dBQDpf6S6IUG7Es2F3phbkWSRUWo+6Ske1kA60Ri0oT2v8C/H
dxlLxnxtuz+P+ThOWlu5A8Wm2dOAQ5wrXPGsL06oAjik7/SC2K0Cj8cTcd8MBFQ+sgP7PD+wy1Db
CTdQmaJBJq2mqSHDXscUee+qTZR8wwNYidS9u5Uy/GHfHbADV4uumowg3oWK+n70YgHr+UMq45t4
Zu6Wu/1IYbc2QZi8ka5gEytAPTN0X9pqIPl1n7l3sCn67KMAA3W6zGGKJ1AjvG1PE3g1CFbxCJcH
BKXv25mGgeKcdz9x3EJELduG5+8tkxOH2Qah4P2oDkVwzrMuQAUqlh0r5PBNYPjcxfANlyaaI//M
a/C90o0skyHB5S77lb0oybeHMJH8nKbPt3DxO2J3aDluTWSSRhW7Cj26U3zTHPSvFSUpcOhYJ9xr
1Y5S+bqvm+AsKm8eQNhj8yn9rZQivbXSvBr40fAWwLqDCZyE/TNzGNI6igRL52uRQfQLMPX7XwO0
J/JuPgjUYC4/eqQJLSEY8WfiB2wCz/Z9IJuTUthZWsUfK6bbb7qy7z7Cr2tfPPLgyXjPFUgDEMan
f6vxkWMDRjBHTae1OBJGH+CKuDQbC7+Awa5B1MTz5bBBDpJukbcmNHZrD8nEpQOSFGPH8+aDpofX
iLBmtfmsMMOPbCqjTLLiiNFixhMhGjmEUFFxTLGQrVEzRvyuJ9JoXUcQy/DaqS6Cv+Fix1BFWLR8
bsT/GoUeab3HRnoIesqnIC5Rb6pTiDvAUwps2FUgXri0U8IVNk7s7h5XqOrZI+qEoPD7Bibv+HuY
VxDNKViaxpywUl68lik9Uxy0nhkcl3IVafm9MunroNx/Gw+L20CMGi9XewsQvnI6W+erUkOI7tSe
cMrvKWYvDFIuGdiungKjf35q8gXDHKInyyPkbCQpBvYqjOduCoy2br/w7dL+DyIyypSbyzKFTdNT
8mVvSbJp+kknTEMqPj7XAXkNpx6IN/vFFUf+EK4VBxGFpba2ANos5LSyVwbJTwt60NLwS4ynjnWc
HOTtyLw+Fk7NWACUeWyWzz7EByeM7sLGoBaJBxAQylpcuHjgRLEzWPH++DHzAK6N/XMuu/Cnkjde
UzNTwxiaH+g5eyTIPCr9VWp7dAUyCauG/zq1132OhaKIRU6JH7VG8mf2d6zjGtITbZXhWsKaQgrX
2vAKgCb7gPGv7ijVZDW4HIjV6ADxpv8QJFSz6rgJfjrYMkRTpJO40JPjtymmgEgnQAeP95pUwScn
lEqo0ZwtILV6eYgM8imLvPy3kR3NUDbtc0IhSSeGS5biufVLSRnxmhnGnwwrR8tM40NZVBp3DIfn
koIQOXqo5xVFSlnHnYrBs8w1U9RuunvUEaT6jHk0ii1E0128E0JYZLMGHwywpbGsgKwu5CFqJPHI
O99+5p3Yhc1okNofFQEXYxWEZJ95tRDSU3gMkVvRDdnxVb+rzWgqBO+Q3TW3xNXXquYwjRnIxmI+
cuXWUDnj/c8p8VjLboTh3lrUkZ6wmOE4W8xvWXtmK7E1YT6Pun/LYxNC67QhENe+UNyKFbkfWUJV
Ris20BgGAnYiP7/BRadeqEo0RvSVOxSfzKeib9c2hiQlbPsPbDM2E/412j8ndbQRxmdSqllOTdLp
EUorc66AVVDt9s/HOF/cPQcOgLyFAecoVzUYf+a10O1NlyDdkElGL0lUqRwtWefTQEv8/6P9Rzjv
5BeHE9B8NqCUudXlq8OB712tmr/ayVDw1wM9De3TCEMEBbAzJqxM0kq3U098zXN2uQi10li5O4K7
55i0zN7a8hj2P5QI5y2wQiAygDfdWo2KCr1tDT/m8io0jbHYi6OhApz7KYlpuO5pWw63/951kerB
mBFYt0LD96UpVUUBWua4y5IHe/Qj9VVoagPHcFECEXJLAKfkI5OYYBYbXXpN2kDqsUVh9gEsrt7Y
pJwqspn/7mpSqY/1ukUvmtMkqtmpIWnhAXwdsuY7AirRpixmsDenbpGVILjPSDB6md5MlsdkAgIU
7Qlla/toUniJCld9O68U3YjCkAsHRT2Gx5WQk1cQjQHeTHiSr8k2XsER509dv8eGDy79EW8y+kZ+
zPXpTE3GYYtyZXtU3E5kw56NETBxklB6/MtmZnnAAJn/oecPwMEVU4gHOBrOq/Pi/KrL8sLw0c1f
kCzkMaZV4xuv29sFuHAwusc2d/kmSTGMvnmfVvFOH6EiV4JrnsRbpiIM3llQxozBdffZPsTpHZHU
DNdHSCxR8I/nuwfNE9By39uhHJOExLMVb/EFJUlhPj0NbpYy5s34+7OpSxEJZM8PpUgALz+jbgdh
nASrbjwbf36YC0QDjdiIp3EwDRA7UwiZcxog76+a+l0qZui4UtSzoJjPUApSUozadXcrqgdmzbKz
9d+7eXWz/EMr2ESfGE5p7U2+FysXD6+/ACOiY6l/F8NgDvHUCJcGlGzA+nRI7n4K/CGlmi3gk4bD
DiUw0KKGm5Nadp6BVaGifdmxtS/IwaYS5oWkCb4D+BLdGGswT6a+NAqJTC9zf/ZAA/3TnlXB/xKZ
HDEjHt//SXVxKF5VEeuoNUFTcwwtOIWLaiIHA4JEImKTJlJjMyd6ZJ2N0y3yuu1YkOraiYNKNSOo
2S0Wolp8QQt/pRv89tVv9m6ZCezESMdnGTZj6K162Koiln6Io5W4dZIoi8qhkekP469mT88RMpYx
eXhxpXkiysD+obBM3G/y9vjapN4+qeIodLkEvRcv36/ZcYZKbNbn4aMFDH53QrlUfSlEnGgfLaoD
7zT8ZgnVvOdtSygeLMfjLFIxsKAdr1rt825PN5H9eHoLk48kzwCiVBq1okIQoUTUWb54mqhFKEoW
nOM+/HL9nzqxEUzeDZLqfVkNFkTLTy9xfq9OWYIQpm4cM57n5o9ovo62XEZ1HzvTsxojzhiT49eq
x7lVHISoBZtE/DYpxtdbPqEQKJnkJ8BsagH/4Vo+1Km9BI6+qRpL/EQp2Lhqqg1La6YCP5J3Le9V
w7VjBxqbVUCYF2QDZZUWGYEue/FLu8K0YK19XylaF+bEZFhogveBPdjUY4gVZEj0wB++Gvs2Fr4J
8BhG8qU9YA4FBesSnxoaxk3oOOhcN3qMyN7qhaI0XWg4od54llBMg1cQCyczUOzDdrOV5jqxad7w
DKNVc4x/hxsxvsyfTCtrEbrcDptIeRzX7NJZsjPujGQCOxeQG1K/7ebWJAX53ge8kG/xnYKfoPX3
3VmKK4/z7BnJfKvS/LKQsch03De1e/ERJC21uYrNYOv7QQ/weil49upmhqnSzu3/mG3zvjtXZddU
eSFSu/lUVVXrKP2VvEehrEDVtTuXk4i/ty5wZDk7V2qlxzvOhft2vkJF2KRFc3Ck6Bt03sk6MTg8
rSMJJh5N6j+e53IP6023hx/IXA6Jg7li4KOqQeh9hGKRs7ut/2fV3A7r4J/BCl+zMI4fY7ZjUAPw
XRu8G3a8yJOG3F7qsEGpMx6cSlTDdNgdEW58T3JhkXflUJXZLeQ306mHt4qPzAygXkx8fAJaO/F8
Sf6nmVI/N7It1v6z+N+HASfYBGLf/hGD5Ay1XbI6g3Y7UzO4kGMBah+2LUOKxFErxZDGWr1LYpZp
AxvbpQaIdHO6XJsxkk3Mx2sDbrImf8eov7Vxy/RHJpPxdRDAET/tNLsCsV4qH6wkb/rRzDji0ddu
DV3VJ3OrqvGb7WMZN026IfcDxML6kX/GZdwYdX91mwQAvdUpWlnniWsDMI6u0jUuXfEwfpcOymGQ
vFc1y60ge1hIqj/uJBsWn21ud8oIVq9EqnmeaqZOCq/4e03L/XAiznPGTE5tIw5/jeWT9hSfdx79
TQR04HaYamaG8rzQoT+6WWXw7Z5eTntdh7qHSpyyDANogFX6LKK8nGf4apTew4XBSqojOmPVRtrq
ZC6BOIa+MvvydV/V+7PVhSMJXJ+FPT1ieelJktnC3sijRyxSrx3sTgPXmYVPk2VlgEo85LsO/lLC
cxhX/DV47aEVSyNFcODjvtMuX+Ku/5L04sDu2ze0NhT+MdItcWAzCxaca8svWJ5AO3Ekp12Dht2N
yubRvdgiPXWVK6p4jMWgmoO8c7QHX+GwlMo0nLKoWDsp5ZNTnkhM0/Q/nAmg3HRM52w5dya3A4iY
iFisjUmLq3kUP4HOSZWdtFVUwcepFOQMAp7Rtr8LXy1Cv1AlhO/joxoe9O/wJxf9B0Bbd01lHsII
YPHMsz4v8S6KUvc6tmfQ7lVftXogE5dm/zlTcxMzfzPytEalmZ8zQBvWA16wAU+4JP097BQzamMx
Bc+fZ4hLeD8v0UFZAr0KtKcd7oP/NIj4A+vBncXs/7u2RgDYmyl2ndf5kPr6vBID3oMJxSRWkOiV
m9f8eRW+WShZOy0pMzG3Q5dqMWxTPKMW0ynZhouuJ5bAdme1JUUM/0fqPcER8Iy8ERtSsHnAiUNA
IuWW1RqXUqhuJ795C5x9ruy6VRJutXJ1utDjhgzENCD7R3N9HCilsQ2Kvk4q0BJnv0gLe2NjkVGx
NztNml5JiinNDcXXROXIToWYJc5RdObmAaaPAAHu1duH7D68e7kg6ZI0nFV4Thde84ful2W9vnRy
+G8/gI8cYdDWcbvHrKag4GP+oMhhA1qbt1es4c0hGMgda0qUuL1p43NLevODRxqZMgp8Lzlpiw54
rmbbDtC2rEodjsKg/aDJ7ridu2tWtQbg/gn11rssSgZFvn8AQ9YqiPfIEnXeFDMmOhRx6gOcFAmu
1IeFgOt878kn01McqFhRx8wllUe81fMRsZuhyrYeV/g6R5HkDEVy3VHlmo5sFdK2k4zcYf4ZGa/l
jCmqv01si5dxtGWuDsMvsVqsfQ4d1q+9nLisatWP0FgIR0D6aPVgOz+IMBHNMUKixygsOCQ7/z/q
lm0lTFS3WbQrhQTkH4Lh9PoL4Y77lzWgWD5bU7NU/uwnr1cTdo5O4MCFM1A8F3xiAUJ1u8w0uQd7
5xzCNrXnrMjPlCmu/9pocKp9OEGJhNZyvPwQPTHpGidp6q5SJv3opMjwBKp5GEvBeo63vD213BoF
WQrsoAZLwL4EAfSeVEjSyd8jxrAcv7CHRaSKLwCVLlqyOCyVSfM3e3WSQChdr+ZUQNmmYo/s6Via
nl4aL/ZyShI4oUbIWG6PKs0BXT2c+hcV2uXcTb+uCPstXvq4CjLTqZTmA9d9FF5jnHHI2KHfKqdn
cUy8QqOqFv0HB838RyeDzimwhNAWYxd0zWgJkUL4w344Q+jKOe38hDtx1jaPjvam4fuzMnOnjWO4
ptVDKhqNWQUvc0Hsb2tfVJMTed11LQ5hLznbJJlsDmlHXIPijCHo1RciVIWAQgF+zpm9SoRDUJdr
tAX0J5QLIJMgHPvwJkQDfZaNt6H9kTWuBUjMgJjtCdUiW/6OpBXy3d4Q1tqNdGybbSxuuDUTIbKV
c5dHqtk9956TH4nhxgd2pLimvIOlZYosN8UQjJD//5KujSkXbTTl98FatpsuUde6YR04JEtH3LX5
fZbFpRtPgGnigwN5S9y2C4ShMzWFC8TWkYcQ3ah10va7x6nWbiFEe6nciN3hfxD6e61ZR8ZWa4lE
YAtIntuKtUdFyOHOGj8c6PfokieigFRzu04zfT3t+TDiVr/nJAE8gdnouyw1HplQSsXvBOl1z3kh
igmf0eK6sKvZ3WO3Fx9U+MTJlqlRjvsVc/1twY+BGSVSARrMn9UfRzuJbJQTJYQUzxie/Pk4clHW
q8W2q65v/l75J9IBsEZ3gr9CIsGXJmg/YzOKNu4uPuSnsTNo6uDgBa4XpM8PmrsoBzJOG4CeVMiG
OTMkAvBmW0Dd+y1DC7JCHM+r5CvzeJ7wwWy12piY+05UKSW31zIvrkT2tCd3Bjivzyo+qAt02Sr0
Wt2gQ0gQ02zu5jly5OXPx3j31+72V8RNOIe9Qdwehhlly9T4fwDtZHcxjk4S9xu5QkmQoWSqzkTT
40p71ueQ1DRSzYk84PLtxrzsdaXwRNGEXUMB2QjWSZH2tWR6YP1ZhTS2NEoXt9piJ2QZmrsRfSeJ
uJfn5+RYs2qvY2cORRafk9UxpPdhZgnNnlSJHEAHlDY/QMJNnFlai76HTsk2254C1VBaSjnQdKPy
pS2yYcxykcz8iCswcJ6lWQUrUHeT9wn59MzDopXaTfYeTmVjlUzj9cj0zAJFGr829J7yuZfJR2L6
TfE9tc1vslIEcyiTtYRltbtEsAvn6lITkGgUH8iOLwCjeRyWaF7KO5L3fF5flZqgeALWoAu/hLUw
nqa6O/A5laF1lQy2HwrBb29y7zIInHHgrdHLx842CajzbVyDZUIVdw0wSZ50nV++xMvpOdIp0Z/f
kTQA8qk5kKiIGhpSOlVoU/5rJJtIF3JPSJ7w9LeBwcLq+QNYCZ/43uWLXNVCPEhInvl47MAQhik7
di8JZKZNqNzsoIJNyIaPdWk4/MBO+9Hs08zmzYuAjDN+yax72yveb+CpvvbDgkXLpIoD26EfMsmD
eV6tOUUT7yQ8kTUZZ2XSPmB49W6rddX+bUG/Vg2BIv+JzdSb0OE92/XyjWqyn7NBssodsO5oUTwx
Qnbx4y1QPaD+1L1/x/ekoKXLu32WFhF9CX+gQbTmbqxThStCBUvZuvu1E4q1NYJHkNWaI2Ks44ny
/SzC2IzdRvQSoMUwD6ACJwWEIiC682MnpI8Ehalpq/T4PolgDVraxynnBH2GNJ1QgMOX2RkyIUtc
KbwDkCAlRc9XvutkogBSkvWuuMU+hVjWvWWNA/yNvt8KVhXARV1bVoRervUlidkEzNrRHFKcbjVX
w+9u43wGXuTdrpKLs3Cx2750geFyf0eJuecKD45i2hnfig8NpAwEO4kuBaX1swtKDyYVJBXQGdas
Gcm4IOxeF1x2V4uZUaLT9c1eHV2/iFqTfrtN2mESCaCekmImLUkAIsP86B3OSSgSnpNCCBobHOLS
Pyq1z0L2vDeb391LdAR+TVtnlNZl4DNnShCdyxVttxhY5UmKUOY9tFghRr029sf25X5slaPdAjUP
rK4LraWmpq0Zc942JdVeVH/yLru8nzJ39MenVg0fo/I5mkE7QalxJehPBXj9gILdAz/ylzFs8MZt
obf00sG6+7BqPCO/YeZLphQf89nXSh2g1y/Yg0sBhrh5JQSYsvl7i34pj3+Y2UtSyRVoa2QRpcoI
o37J/o0Ls4y44WWIHs1YWRpQx24ATlgJe7GYVIl9k5InaGKhHbcRThanaGfzbt1fj9bfzwwy+KZW
gmBxTHaOo/GzphrQ7HofO7KwH9kiEkkzO5Byi5NBVxhMnVb04BQLf7W7Ed28hVyMs/4SbWHVU3kM
Z1UZXnT+n2r9fyOZ450j4MP/5z1WUL6wyjq1h8xOoS5x7jj+p4xVxm5I0GubHsU9VwxdQk5gd+wL
x1Msml3cf8MYZnNarSK2Ajx2zvCcxgsCacMn8GBNdqOpXpb9i+cPqV7snqip0GEsxWyRPndKhx4t
DNW3ynMrTX7TJgKenlt6Od4Rb37Yg3e94fHWAKx00mYpSgoElYjyRRjp7ziAixdPgAXds2ROyPwf
H+kj8tEoZRo/QbTaJjSOfouSwZiocAYFWf4Tm4bgpTiFeMpuVP0HqjfMas8Wd2H+E+8f6J0tJ1/U
SYXb+Gh1qhM8j6mDSFgfpqJ3UbP01xuVz5F+wzJKAKJL3sBluJeKR9VDVjE0NthYY84unwC5NKhk
skKNOKMtrkKC9WzD+StKJFoXGcWAusxKG287DulfcXkby5g+i+PJZka0lzWMcY8/uBLgAncKiuuq
SmA5+5hWQ4a6JUBvrVite68WQ3P3T8GROjLPJBoVWcrym+iPcMRA515p/OGtLnFHWtT7wA99VRY+
qaNOmvl+CY+LoQAG4RbwiqraM1Na/nxkSKSx7WSNgM9vEObUIuK+LEKpICV9PGKVD+glSJTE3HwA
sgYxSd0KWwK1kP5NJCJSamyUen027jg2xqfzyCyeMx+joxhD7g0J70TW1LjixdRfZkFc/GU1moMa
kCcAUfJRtS66uw/jKLHQSwvBVDUAXmFyChLPLQTfv09YShravVpuMcY2SEH7w+MMSPrXI+W31kq3
XrFICQdCG0/PTYhB67v8SdWPNWMPnbX0zk86Vw086/2Osja/Br6h/MSw6phdbwc1+To2TjkuiFMy
rj6t5GgeqJ7SxjC4I5oY8xyHe78UvqoFe8VEBVNfisgMmqpR0VJ+PadoDIoskzDP4FOKeMwwOQyD
fnf81YfWsZJfm+fGn6qYm3I+wSsSIPqh00w+dB/H2juX7hM1QCysrAqveeWkrQRDBsLRcjE7//X4
H5anamx/FGI+SDTu8T+9+bFeKL4Upd3nm3AGorh0JDPnMixMxZyA7WeoQTLsOniZ5mXUTmfCJlC0
drY3Wa6gbQyUlJ17Uea91UgNZK2HB5ZXgpUz33zIryRAFGIiqWtZP20ysX9eZ8kusyzqRIe3D2Vb
050+8lGqJXzbN5a//VVcZ3UB2o5LBY6fH9gb0kgEm5pcE5Ydue4lT26Xf7OACRwyJgexKZhnQTA0
sjRl8if6EqvqebPzcY2k1E9vCG8Wm/+H0kTXwzdshmPtcCaLLLdGIavLqhQON++6fyNjkHEoWxDw
QHTiZlfixF2nZ1in6RZsn1nQ7Dq2UA7DFvnnLDoGddLfm0ldV9q7Uda0mYystkXkYlaEdsj5Pukp
629oBM8X4psx9i/Sr6PSSCQmDqfEUV63RVKdeMn2dA2/cNj19wZ3tOg4/mzyMQ8FLL+nQKM8DslV
tjj7k0Q/CYvHxN3KD4kfiezSKJARxEJzD5ekMrECFKcrEsEdTmOXvwH3kGKKh7iixlYJhaDt8K3q
y0zmbPi5RTj6JjhB2Op5mmH/tYuRqy3EQV2A7mELa1vnKCDLW0YDRQp+oCz0I+EKTN/RFX+RwTR8
tyGtJFLOON52GnyaAeDY7/u+Sd8N3iAizrUHdxdX7VP9at8v0XkHmDcr01jyW0c4plZhphBkWbgm
rip0GYMDlEzcM/NAabs0OBtHWtMIiVVR3e4lc2JOG9H0TGw6UR/GDaldJTRMoQD4xrjaYCgW2AYv
QjNFof7jrHTuakCrJUic7f6uD7Kug2BQn+PjE/lx1ms+GBkXdKdgpIoTLvWyVySjxZ+2k6Sy4yWd
F+qSyDdf7nKp0XiAqxuNv95OdXZnR8TralZPFaHnJ7AvDYpxRKS4EU14Sk1InfTh6QgJDdkeLzQH
RGUznCfTaWAlIH3zeEt4RzuW8AJX6fzZZSf4J7iBUWwhM8jp7j/Dw6vFtuZ3s12GQn7FgAimjVtV
V2gGX2wYgj9svBCGJT6xQ49QBXzOpUIMbhUWnuhNBnx0advvcCV6sd1BVX3xy8Y3K2mJe3YUUb10
N15kTASUOYhjzbIBGkbeqcoKaF1IVr2VSznllfIKAPYWqHIfQV9y4cuMxL9+3l99eNaqo84fcPWj
bm2VJmBcgIHu/NjxlXb66rEVPncF3dsnvmTAP2vbsdDecv44/phwaGsoQ+OhGvDk3qBBrhsTVKpe
ECbt6Tor5joMDhdLi/3E4y/AfBDsSc5gu0fPIA1OtIa9CRp6DgmrqmVlk1/mv+2ec/0y4ApDRRXp
O6LKK4ZY+aOoO5Y1UGPUmn0SK6FIAFN0C9mMwmdq7bfO9gXdEv45ynzmQaCPbqEVHClBHMGCpz9+
Pwjrvh5vbb9P7QncHOsXIR87OhMSVvbjJXf3Jiicp8HDJRHpLe+yv4vzIvuw51zdA1JHhDateL3K
6nOgdONy3C69/ltbkdijdcT3/7/JsejtOqorwjLkvzDrDF5N9UZpyG7ZOQkGhJ8qT6qeR9N0ZuW/
KMPoHFsyCqP+4jNb7xT0aymxuZjhSgI9kHRXpfahPfjxPrJCymD9ITccqZ3F/vPOkMFFu1R7GvLi
Dbw6QpiCpB5p6XctT0A66itDRuFCKm2zB70vMHJkpnR0VhC1mUNTwH4tqkNUMPS9oYBdcuK7nUXR
EZ36CeqxYFbsYgMQX+XKfoidi3r6wIiGbYrwLgVp3Rp6OVAl4U3j0Ijlng63mHy+UL0jF3OFYhS0
s/n7YW726/NDU9aEEzlzbCYQC02B9wiE5x4XJIfLMWLJhaYJPPgHLBLwi+7h6LTNlcIkag0tZG+Q
P/APSwTM1oOWNkGghqJmwwcCzZirIYjeJ51Iv6sg/3u2qmxVNuOG78+bT7lmdgVlmrmkbdOYukpp
ZaiRZMLIiBxIr0Ezt1HtyKb7qNg8VkPm5Mih3oT6Aq7M5yoZ4eIjd4CsMIUpOevzxzG7pzw0kU+p
cpUVwUL14/c//Jly/2ZmjFhEvZR9lu06MH9Z0ZfBNXSKYlRxA5hWc/RfY07pWbFfpfa05QaCo/uM
/O6mGE0qPyIfuHN4oPjYh17FnQC5zomZgKhqoV1bKBW9/y+xwiZyqZzy+PoofLcxFvYpWrCSKFnS
LNNJTi3/+PupkBQnEH6WXFyvQh/wuGU8RciVnTH8IdSR8FSzg2ChdM2HD69lv/YG0Y9cfKposSFj
kDUwPkk2HJV2UHEI/0+vqv/kduK03DmbWgATlLKkVgb4t7LVyZFjHswmEB+2tX7ofMyredVArihX
FZx7KcoFDQ856/qXBPDyGZ0Sd4lIJy0pkyEu+7lFo2jDF+cF82h5Vky7aYLnIlzXQYpddktZ2BLD
qwvvbpwI53PBcMX6JqqlBterSb9m0x9mgGEnx0Ld9o+4jKqhpc5qqTtWz15GuocJ2BoBbKlMtJhC
jEODrq5V9p4SsXi6ClGuJHswvsDINJvEXo6jk+98RcNIwzXuxsjoNAKB4Jv46JsSl1ByIXreA10U
QYAyoTsy/qFLPzsO5Sp+36inzGTvgmPQ6+80HEZxzl28IhLBNdHL4UXgDkC4vOuytCqiJGKOxmZD
EoLDo6gi8Ip9P1sawBQ5temDTTbUbLjRUV5YN1CR9Z/PwENeaVllsCeOv0VmitPt7brSorosm2la
RK6D6vFjfyouzxj6pOOacPFS2Uwlfi7N1otYSyrsylCdud++y/7hAncQlqZd2fnPJFmv8oI/gJgZ
H3D/Z30DJoHEOoDfw6jxtWhzpsCmVBgS0CAvwWmvNAIIV2BzMd7GeizwZoknGiBxTqcRaJdAIqWq
GEHUoOuL3lDG/F67ty1TT839clnCvQ+hb4JqBlXojCcjNoeinU+7BZU5+bdyGh4lmSLYBM/42cih
FSo/mlerx/eVR4hQiQoaVMpFoVryk529u/osFVwoh3V/73/b7UaWoWKCicvT3fYia8YygvZapUg2
qZIAR1eEFz5bKdDs+pY/BNcYJl/NAbyTYfoMfltcW3w9lWDUvyQmD3N5q6p4wU8yRjctwf9JS6S6
Gde8V2YmdclWFNInBXZWiSS+YaTVV3AfdRB4BLfPUpvRiDUlC3vsyJH2ebL5Ulb6jkUwuEpGgL87
g2qidXQRWmpF7gxtcopRl/zliK1xGh1vqRaic4JvMk2d/+l0W5ros2p+NER+E0ev6aHhoiyeAQ+C
q+HvJ/+SG4QAlAgsiA8D/CVza/cOqkI7H4w1mXGJmDiv+HADWAMprgQtoVINJcIb+iskTPwOCKAq
yR76tJJHATLeJPR+AEBp+65Lo1/YAJlu8xgkNaqXiXjfaK/XAokzb/FASn0uwurK9tlASPEwFYDr
sroGplf4EEIzmOGYVuRCP1cf8dRO6den2HC5S0Z+nzP1g3bWGSLrRlOQCKf2WF+aJBeqwS8l1Hj/
O7K8cFSx6VnMAcTcHU6T+lV00JRxBFzxbJND+mhO56/pFtRxOuaWTwecUOXxP6Lt6JZPJdqpOsOb
cij8CWXkEqZT5Mis3SzTMeRog58KziCNGVkjVbzGyTnITF4EGat9cwP9+/m3tV7f5aKZblOZMFKC
vo9j2W0U2ehiLngM1CCkHXfXkzhDlMixHKUCXC2KQ4DLAfXl8oFk5fPlySaEbr2MdJKYvNGbg2bz
ZawQHfAm3fp9PkKxKCVWjQxn+uHEAoYrZPQvvcVkvt8Z2Loe4P7XnLEFt3MBgVRQZIMSpLTLyv3o
VtUCTK+kWlCHQBm7cGHTY1DkZvYVtIC7WjHoGEyka3GHHRb4vgsO91W+GdOSJeS0jXkO7PmRSUGf
vBptb2YfcD2Jvpj9gsGSW+4p8E3U0Sqfz21wwyJHZrv5z7Jn18UX973QMCx5uBQenrMPNXaIHIKb
GZJnjodXkHgavwZDZ0pArbdhfBmS/Sqh1E2dRAnjpF6rQwKmphH737zsGxY+Z2N7zBZGDLtxsG/L
8l9L4Ui8nHnJmAlcWlnfQVUB8o8I+qGJ7ID9ppd5okkscAW8jJiJ5gMfqudH0Dx7YSG/Ch97uvtw
08O+fHk48hhx+lsVMFtOaUTGLHk7SBU9lH0nfT1eXK86McMTiwqnwwV5jMYoB9CTCqq3PGzdNwBg
peR6e0O6yjzdd7O+xobgCubhpbw4Gq52xS+OQarA0PR/jw7TEEZmxIxmi2Ns0hdy2Vv1KP0TEf05
0q3ydtyMSiYajuCG3f2937FKzMLQ50wcjEu54A8rn/n0Q+gyiZxuNiYPV9T77qP4948dCJhdIzxd
TtLIXve8AY0d3jZSYKJiQUtrCjEyMROp779sUjPhOrmv184WYn4MAUg/xcX7WtACRRk/11y4ErGQ
mZv1DS8i4r+Pxyfs7VpRahkOyABK1hu0bjqAePN/0hX5AuLDiMykkfu/3oud/zfOH3PNw/VFiV7K
rvR1mQRcDV52hprAEsT/DlQWNErlvF2jgc+i9jWo03HXjwuarU8pvvIbZxH2Qhxz/RTuqgso1XBC
BsBKrwBSFLwKzD8eMMZ5p3UIl9UB7PDMdzeaNLvKZJorprxWVXs+55i0xB1+q1ShE5hlfm9YIoWi
Ny8slVRdUM55hE6aePTc02SS0ap0TLIP9uFoQBUCRGbEuUuUDr4ZX4xtuW4OJ19vvMlYGFeQXpES
W9tfo2UgUU3dQBM/T3/h4pXIvTh46a0uxL5zRurZnvuTNyr0xlbrQb4ITJ38ofCMIbD+w2APbrHa
whSFYTvFSp3/+r8XhHOuslcBeDZgyFgJnT8QdmlW6jgM1Cy4CbmpZVYFLv7WQVbKfkFd5tqclSmH
PsjS0rmSFAv2lYiknnt5/slvLPRSBVt25TXRf1BNKa8fC8GhRc/pIkfOtA3Hd682yVkutuQEBYYJ
vWZJAcCTYdiPqj3A3gkhLyn9SlA5W0Z9Ri/lbwwehzNOKajW3zoksSLbc5A79rSyiVP2UKwWGqf1
QiW23cLCeBui9Hrsp5q5ivsCug/cnaB1uXfwdJRPltsus8g0LO5nduB8ff03lC2C8hm8GtYqb9Wp
qYgR7roVxCJoUZHTNAXKjZBLhfOOO6kUruM04e28VmpBOpOZu6vQDnPABn9HFMm9J6zjKuUoHFdT
2hMwAGvncyVgAfhfksPVwzXI3iI05mytQHWypSJ34Zq+GbaeUkbNsBsHeqhzAJ2JwW9Ex9GT6bhv
ARTSiQQ0P23zhgODuVFC4Hn1jU2JikdfYbOzmh0144mywgf9RqWkIt98g60L+GX/XJbZhDfyKSuk
FzRdJbcw7bM/2s3f1B9XEXRHcuhNpUftpjhibt2Nf/y8CGWIm20NAff5NX45Olj4fZKSrHEZJka0
M9rouUyoD+65WbIOW8zOGVgyscvbBYofXX640ck5/XvV4VF+olIc+FN2d8T11oxVs/+ULn8/lPam
Y6ujIrKUCzMj3cX3lrp8KsMhPUl06VTVnIRAweAU87koIJJ6+DN5t0o3eNzFC5tsdqs2zeBCUKk+
BwUuVIvVcz3xUo60U+rwyoB3ZtrFuHyvLN9NyxvweEBQk3TX3sueeHT2bPetL1xuTODnuPtQK3J9
Cif689WCzH3Ojvv12yQ0PZTub/A8VRyDvG9MRmZjg91ClXGBjG7OxopSHFjH+unW/11V4+fECo/E
ImUHgG4haz+JSz6E0Rt4j0I5dM4e53W7jAwVpdts2W8mVghy78emdQl8VaJauOqLFxFgHREOhybH
VjDuhl5fF8q67BG9JkJm5reTOT8IkE4Ew/F+GVW8eePPG7MfqK/+88Ad8K619fhWkC4rJArHALvH
1bDaF9Re9bFFbpf1mnCyoyjXNxvq6k2a4YLUgl+tc4GAkVMFZZCg9Iz6UJW40QOhvdILocFYnXXz
T/P0Wx/dIedhUU+zgiBBLZcJZ+rLvb+XFgF+r6actaMEMuRVRluKo5S+jK1z2FrN6J7FFzxrqsNi
+PunZlOesBv0P8ASquzAVoX29fQifU+2FrxAKCxl/OzjO4PAXox7KogljDnIlN4/L+siygFaGMAC
g+iprttPyoQnvY/UPTRXT/yK/VlwE3iHPoSGrNV017mzSymji9y1NKnDHyX3hP7KsXXJDRXDpz5m
WxNyKymhpK9+sgk1mb9LYIJ0TRt97aRIFYTKOxCL8diwu8Cj3//nz1fF33VruNtbhtdbwj3OG3Yp
mhtIh2mNydqjuY8lzfaAApt1aVGCpe30H0PfXEdGuowBPDECOZ+j46+mCRR6UmEwnhlSQZAmDeUR
f0wAazxrbl2JiAaSqQ0JyZHbaa+5fpi/h0NLfCMA484hBDcJsv1hSywMNmbGdb6eO2GNCmzlZFs7
f4q3/xQl3LcfGtlp88Fw4jxBMlyBRQWND4nK9JZBUiDzWFlG2CBIUVDAvC2OtwZfHdUyzqP2d/8n
nnlsKDjMXt9Ialj256xObuV9mLIFmiuj7F13YqKZrAr2YZrXfEdp6J/q519E2HQ5hHpFglmziXi6
1WqxFmiEKSx3mN2O5oIWcQvGZuedF9SPx4r6e2ebWgfClZjJW1cpOAvctLLSTWrMNpZutZgIySec
gsuGn9JsjKWVfjAjDHtgZfCTO30fKJlPhzKvpYVbwhuUXXbLDpo4mDxEUGZ8d7TYQCkdNs8sGWhr
AFuDr/TnQPRDMHkKIIVG4owvkpzmACs0wwRDUzQYDGDZy8O87GEmL31Rii9ckOF470eGol2DcTDk
InA/yrEEk+N1MEH2RsW5VwdRt1/zGGC4nHT8MdpRM8D8a3RbiEQ0e0bILsiVmdLrIytFSOJE6xDb
hNf4gLU3OfqQ0XuNqCbX+8L4e5jrrUc96DFISWo3MCKy9aRCEm4J9BZqX147He7rCAW+C6pg2svA
qk5oIoaN79/BCBw7KR+nH2RuL5Fk7zjtEXM+LQTd8bDPAhLgHGhfH5H0lJQXgpLR2uWgoouTzuGc
f/C4EACE8jX9tsD/KOS2YepFfQQGbM1LaNxiIGRxcA2KViuuCb/rk/FUgGRorqKJozhsGe6DC0mG
4T0ca7EzGTj/oZ0ImC30p0N4zqKcue5HJ0lOAQTKWRelJNx6UDkZDt++0ywjP9xjYfXqUY4uNvOj
56B8UoAuUwv7xQ6+0le/hUxgK6q6VOYlM40g4SQCxzVZBI9YEOWnU2hBu+nPFIKUsu/lmxqg2J/6
hOgNQRmB1/5vOGb29mQ6qZWLmIMwy9y/UyHVTnEXd7vDzjw8jQ0gUllxP/hrrrhHf6UmpjekS55f
wZuxT/wVOLzLVHNfT7QkX9djoVeQ0fbr8ZRkiPwj/c1T9sdL8e5AumYVtUHOLwilaAknoSROoLjq
7ctqt799dEel5RiBkAK/HSCASNtkfPc4n6ooT//JDxt66zPIuArXgGEMW8WNcqcrLky5J6rFE+Tc
IukG0LVkGhJyKxjCiNqHNf8ii9OX/FeOzFFvE5VoBFRTMZq9QaG895e124zW75jeoOmbK2dChp/1
K7W2yQXpqyoEJ+c/Pb2L/1FcqZ6Yvh+w3SwzSPJ1Np5oK70YY1i+tl7Tl9XE66nMAonjh29t0A1H
OBgJ6bbK9Fv3k48PUQulBTjyYqvf6D+tfECQTepG0BntjsvmoQRILDm1GRrHY+QuwqjECFEGS08T
8LonKB6KhKlGIGlRcVJHtlMO31PySUaYwFsAZFQ6/1gVH9Glh0aELNaiN4ucyXbJsXRaGKPVR5de
pGazvbOech+9jdeU+fp5q9YAiqRyaf2A/aZJYuxaBhGIAt5C3aJ6vcmyc2uRhoVEz9A9f8MAE0jp
wH5ovjYjOhcuPDFzwPl8e7+T6jzcAqu+TMMDkmj7cDvarEWAS1x0NA7roK3IhuQ9rv4x6hwZ4HQp
7MyOPM/IhN3WFyVu6+QVWuX9JeiDyAveH4PHeSDIB9G/qRsk9uBchJA7jKUEfQBpu0iQDWP7ORcd
NK+BNirL8kDaUQJewyc9dS0QZyFzJ5MIR5EoE+qH6qwrs3HMCrhYPvFZR659ITnSl1ZSri+Ketfo
o6fmBTccrhdFQBe59yfMYKa2uw06KH3zW4oW2sA0bYsyBk6FBIFDqXWI3AiWWNq3GIUkNvP2cmtZ
PTkiAMYYBYDfc7m7ECL+2KYLRbQRD6zGHBCri/DioH9QkWH/W2SBdYPb976RbvqWU/qRVpQ6p6VL
eax8RS7B9STUqQ9/kZNuY4VRXvUV+EXDGwBZe/YaJoGxhUbUHmhe+ced4jMTOEfsqGUibMyU+G8j
eFoyK95t88fDGKnLBnzgQBpPWzCt+SN7AKirfSbjWUN79G36bJnHV5Rq8Ma5KhEGOAwBmbadIldr
K2pTOGSN7IPpCkI1NSBzoHmHueDojCMBYyzeLm4U7w+7i7mDYy740ZlUobV6jQMSID8hb5CqrQxn
t1kvwicd+BfR6ekt/mcGAaeUaxA2DwgIkwf2Qvubuf39PS7qLUpWoUPGqDwSY1h3QoKvDXHRKKrp
RdXKWX6nAEax3YaeK25QYmjz8vPpn6cQvOyaVDkFUyxLwTsL6ofvrt2FLDi0oK9KBVZ23GQPBnMY
cTK4eipLPaVNzejIKYlGEIe+Uk4/pwuEN8u86W4XngL7QWUcZk5EE1WeUvRtMQsgxQrs7jkOfo2r
F5yPF5abPh4xvC6O6BpKRBiKlKJ2gQXVEdSv1zldL4rLPhG4bvlCKp8Xo29BxdlPYbh/4pthwSoH
WeoHTF+IhzkkLJuSVfPSt+r2bkYjZy4JDhAVWYuPrAkqAAa3G4e4MZjt0aYfQEURVY0iy6bH8La3
OlSZAUSRIL5+XXP43gaznZdUTRgSRqsh6qWujcP8yEjdPCTALYEUWkS59T7t+R6+B5HWZelRbxuJ
oyGVIvQ18bohsnLjjoCNsWVkkry8gf87KISKdPeYjzxujoI6x9L6BW+sHrdc0kYKg/uD211yo4nR
BPtFSmlVuvEXHctwz3/HOm3Bsp7cxUTVf6VzrIcs747bSg73dY6IjtnjbX4bLxzQg2NXffbPu8Rb
9f7kOv8TkUdqddEm0hqwmslehzw53VesbgvxjLIB3YIkCqD8nGgxNW52gLD3W2jIF/lLIgv0a5Y9
SuNbT4s4QxvjaXwDTFyqBJIYgJBlPNdM4DBpDM7h2fuk2K3X3l5Qv7YJIoVhECqoIaIsf5AF3WdB
wzBjqnE7Ixwrzp/djtfE0Q9HZbvgOZDAp326rP5xOCMMa9lxqaH67RDw4EncGIZ9lvXrWEfc8xuC
SdYsyQ0M4fkuKA95gGV02HrIK4aADbyCkYMVEUzl7ndDuhiF/d0mNvpTTWOPSVCUPDz16jlB2I8W
SQV9QG3h1ZSpDMM0mltsEFoiEMVB7grx46IRPnsTE5839BbKpJqMTD9laWM4xeoX/o2Zf1vxHNKW
Y4srZD9WGhJpCaeelGgvKPDYneon652uAVTJMA4sRkr+QK3R/G+mur7lR1sBuy07bIEjRxlDqrf/
j2650cwxoqin6y4CT3RIbGxQtHMW+wnOskf6LOy1wcbrk2zlp+UzL9tL49j7Qzd7sbpw/SqEUFl8
yIXIP6h1hOUMDA6hxKQ+rkdmmLFHpyVZ7R+CKpz46f21JvfxuNw4k9pla5TgKF/s1qwYaB0LGFuC
pXtd8wsQWhyVaLWEvt1ZIBceYWbXAo2WWPw/2jx6P/0l775Aa08JbWXpD555TYLJ1nlQJSzRs7Io
14HMKKqCcz6OUAKziV/dndkzj4EfoWe4/2dE/bffOG9YJ31RqpqHumezUySiBaX5HT4av77GvvzJ
bQp8cDQ9fkQEecmL9XQswFLTFz96425DMkzgr+qPraBJkw6Ldf/vClYrZvxrxwAaTWMMqW7iTP+P
kQ9z2OgeQ5uhDV3JFpMV1jMlxZPc3lH+fak9kO72U541VvBYad5vDwtqLi5Zaj7/Iq4dEn7OAIBK
MVeWu+km3drydQhzZFN+xeIkgrRfCpoZheKUgGLSB+kqhiyaHX6lfZL7kw9AN+6yb9z8pwJFVnvd
7JbEiPj9mqbtUm3KSNsSogg4XdjrR2DgibXhQe1gRKuKg2qk3vFaytui5sEE7Rq7fZpUriYl6FcW
U6UQ89W6pIsgjUbnTixCiN7ROl33oQWVDYLz99EwtsScGGSXrv16/gezi9hLy2xim9mN/iLslySn
VonE2S3RaHxtrHHP/I90qu1hHG8mvArBoMPEMe12/hCI5zNH6RlCS33imWVC6rAe/BghhUqPShp8
s8nVzeOyaPhDGwBPVWCQ+zu89KgvskEjqTJdlWS4dn/zA1oy77lzKogZ7++2I9dk/r+NCcJif+OD
XjlccztuS6tRcTRJiItr0bqfpYjsX8F0+R5fQCAo+MLGUzP7bhY7QggNgmiLo4kFer5hRYR0QBQD
u91m/6GgQQTIJEyMGscFmuBbTuTuZfIYALNc8yQsGcJJTw4kqGaDnctPMMxGcX/j3VaSqD2zqp4L
A/73+JyoaozpHX+rcY5Tlru8KcWqhc8VuqBcSixE4Mu+4ZiUi6VqBaVboYilS4/443oqKuYLJ5Ja
yiR/7ShILI2HJwPc1FuPs9PWZ/ABVjr2Z6UrYCrdYDU4URlf/mu0BpzrR7abRFlAzZW9CM/hciSI
bSCL/TW040XpZBvVe4fd2ZB3cgrbnJejdBFoamJBLPIgWvbsouRnfF0Om1DgWJ3p+bMuHE6x6dx5
c8a2lJ7lTrRbNjI2N9yGVjVlYsqjK38huo5noWrMX5TQYHcDABqtpJxWY5ApTUgUG/KdfclOO4IG
9JQrgTtk6vy5xfk8NxhDS/ONpbHnKHn8xW6AHBgBV3JQm0tVmv4/ewfnAaiR9F9q9V2XBAF79nim
heZZAmrc4YRUghpfiDAb1fYl3qHKFe52ooJxsxsEQca29uj2XLQUmQAMFxkNxo4hAZ3zYdrYRbzX
libZiLE7eCpN44F1wN6/usun7bCjpnN7DzTG6Uxujbg+FjqcHhOAeL8ojmnCxlJ6VvwgNLaHyvYw
IJNKmrHB/zqgM0OLm1yEA9Nw3sk4cF/mUOiqsPlCoJwgpD4j7sut/SqTOGW0hcspUAex2JiIhQ8e
6HHrUJCPDBm7sy+LgvZSnDBf967IujvAWW8HP5xfK784zGpBosMu0N7rO11slww9diIBP8BNMlnR
tvFgMR4AGw8mEuHKrdcCoKuG20W/nUhyuU3d3f8jLb035oDXmPizuFSnG4QnjWyMxFgAx2/N4unU
zKZQ70UnD2loIJ5Mn/rWWhdXZwA1bPG1oCzTdMV6BwAl9zkbwdArEFRAWFtFS9Ew4tKmnGMXzN4K
NBSiIS0uAghBD6FznDKJl2KUOygdPlKRNBiWtC1Eu6uEWd0Ro9c8e4fso6E46tH3WXvVjwQ/cl2a
ARWk/KISQDK6awJVNljiy9YrNVUKVjZXjz1gyrQM/SBehmNtoxt6jmesraKFVYuLR//Gv4eEuCMI
SLgZ9efnaO5zgPcb9IQ0qVMRJjxktjHx31uoKJ9nVg+XVCCJfyn7y0I+3dpEbgbIdd1xp+LT9GQG
/kKey/l6qgf9TfZnFQsIdETIXhLEx+nSCSgibbrVpApnxn0GXdF1Rb0hJwvgRcQyWYE4w1tFkw5t
s21oQofhETQJmIHZwLQbkmIEPYkWrSJnB3I5FE4GZILuKllKO8AGuV81EQl7VNglr9D0ARr+IGMK
IH69OrgidmxgSJ4SDl8rWaEUgOMr5f5dWbDQTmw7Bju5tK7X6p5ZTIyu5TkwV4ukIm5iVW5Wmc5m
z7iPG0nguMmzYS8iJaUPJVa2S9RVjj7YbjsEerjcGZngmhE1/XTiUmbNIxCPz6Qx5Ad2QTmUbhGp
PRZIO0Kd40VppNIkYp1qYEUv29DasKXC050a2rD4lfg+EJdz0qtXoAcKPIPq85We9nqpIJRMQA3q
x3N2SEKbMkyfvKjdWtivFhoBhVIV04vAvjqJxOMiA40yOLURI6u7ot69aUwIX48CS9xPFWdK8RNj
m/pKtyTOWl3F4Dj74JxzRTCOWUhN501DQ5oYN9fZaBZWbZzrZ7hzp125yvGnpq+1itf//Uj6aQ5Z
pMgnes4pAPE21kJObR1vh63IKFZTwcWdosNB2ooDXqG4ZCYnXXI7c66esNYa07e+/44hvyTnd2Q9
Okp/d4hjKXyEM403CFaehq7KD2OM4bjhZ1X4OpFv2zIdy+8NyUemD8RAItv/0tkBN6z0cd5NYiI/
kLDSa9MZwPJ7+ZwYjIzz4xEmNEoK4tu6hR0hPniO4wjROnYMFOYyXRxv0PKHktWZblkDe5VpyI5E
k2CsaQP+99RSVgkX31goinGk6okgcZPMcd2pWsf5JZMBpwjonsQd1/saKUtaFv0M0raSNHD57Oqu
ptvLyTEVIqk48O6cGDohoLZB4jHNCVKGPS9ztWl61XxU8gp60FhpkhzGK8KY/+VfsT7njOCjW4nB
x9zWJ5LXhjJ5An3+uU9CsUBO+f5oVtBWbyvoXg34RQEl2Fpy2r1ESYHYq9KHOlGH/aV5kH8LvwyI
CLZznhDMIQAV0AOtOyGQQD9nK1lmT5MeNHgZtg2MnwC1SxfoYdHmgXnIHjFbGF1N+btsm/g5S4F0
6tK0Xx8WyOri0AOWiDoePQAtC9N4qHEjh79hjm9I5xKYuO66TRlvm7uaHocfDTkT5a+Ced2zgorY
KBPtYTT3gWhW02ENL4IW4D0TC+Kjgx0AuMsspmD4/JW2OiuoVmr+N7BqHyYWOjSgQ4miX7WgcMCF
GT2YbFEySiFlBDf5dq8zaKdwlpzVqTSKIlDXhAcmvQf1BqUdcALi3J7kqOlpfFHwFmU4rYI91E46
S6SZrZjIvMIEifkNjOCIAeYKLV11xX2brobFt/UsLRD+5C7DPtwJGupJygWgTz1ylBKsMH9h6eRF
V91M2ZjqtAUV3oWMe+tfQVRM2OwuczuX6Yip1mlMhpgGUdbpRKv0dZ+wLlhXu6+ixVubaZVb5W+o
Nd4FVV9Y8MXZrB0LqNysPMmjAJ/Y/brEjeIObtX6k92VXHYmELeBnhlHtBgZ8pceyE2vBNpfKlR0
5OovmrjOaDd387OvfqY8UciVaK2yN35YLsU3UnXaJVSNsaIQpfM8pGuc43bJwQuJO4O2jlzZiMPp
bofHmv44yKY1o0fKe2KLWTjZ7QEs5RWnrYezsnKTyCad+YRXEvdjjTt3Ij27+WjdWPxVyRuUb5HY
YGwutN7/7dht6qvLhNklJ18RApkt5mKI/yrRUu/UtIAHruwJ6JnJ2ekIozwadfffTVIPF9FIevPb
oFfWtClRia6SUOpII/JGbt8TVQ5Q3w/U2NMg82W/lDJi5gXMtDf2BEaHhWvomLN7/nM1mGYnwitE
OmRjArRX557sMC6MOnXspTrwlpcOhtiIe3UsweoBlOlsoAOQ/gMmOZWXErGxRNNW/H+czr3vl7gl
6laNMk7Xh+KxUAXEwegYcj1GkHa5wJe6FXYijfKkkKXDRuRBzMUE1pj2Sk2/G3sI/oL4IIq5h8uS
Df6YF2tnsqctViVuGWuaA8GB+xLqzvC9/l2t8+O8pSu0Bg1bIfrmvZlDhjUza5T93t8CXbFYqsL2
TMvHnNUnwYkamZhPcHtUgyM6ipjtNKLtfYb8j9Az3kwpebj0WwLt8Qw9ek3lbT/TqJRqkGiY0kwz
ZW8YPdm4zJM+lJpIQqVgS4PKN3GOaXqwGHBSWyECDYlzdnU8pHdX9FkwRMWWa+vp06bYnuimn2jh
EXiQTSMLpR+bB5B28+3Ux0APNkQolwGOCrf8MA2jT38EFib+9gdi0/N0Quj/DQ5e/pp/CScWFcrn
iUnMlKISlh9kOkUIxd+VCI402V+KOycOw8LMHBQ6UYjFfyLSB/FBpTPCfcdDdw/U+deUYNUw/7O3
/INu1b8G0RdjrvvgH5bIZH0HXp3E6s6XhXbDMi093es/gapYaD6M+zDOUZHxIny5dfdmRX7vgfzs
2dp9cpQmuAwajhKvwAtIR48e9eS4UgT+CHj/ki0eG0g/0iAi1Y2XOF/K27hOfEb1ziyl9i72Ad+H
/Zp+2Q7GXIIvV+uo7u+4nF+EM+WLE9RrW4TfTVc47DyQjC49Fpltb/arcxzypeXHQRhhTcW2OslX
0vwR/KgT7CQ+4mEXd1Q17lBYaclScihH+vbojea5Vm5BGutPj55TVzO3qUIBvxceW3K0iVc1iHIJ
DXfvmgrGgnDkORcS3QMZjOqxaf6GW2ps+JoobUDgSEkj9plwKLs1rmB4WMNtSDoJHQ/GzzmiiE7n
Law0dRzCwwO0hEmYgt29BrVJ+nfLC0DS9jxo5RrFUFh7a71XfAe9MgDyAcIbz36vKhmlrFoHfhLs
HIrG8pzK5KSO9GKq60K88N1M8VPMIQ59k5nPYXwJcIcT0be3RTLZbvpThcycniz7pbw/DstIrqah
t5UfKUUoYx9aWTtNs+uptfA6h89loSL3m9nQmQUOVU/BxFZiRxtjyda1FE4PUYALMVRzXZMWD/gi
J1UfC4ZNPgS1iBV+3lj8sKYjP8psd5mj7SzhuHKtztubJNxcZlitxF1HGzY/DraVoGfk3WAJNMF9
Show+v9tFomBIbGh/LAm/SjRkCCTN4V2c22x3o+EVuhXvDRJ+VZAPSmQsREbM2+RCSLqZyGrEEdE
GGnDKg9mH7iiCFrpkETenmN395B5lwkQjf8s0ZFIKnaG6n46YCszNf9lBZ5EPbrWQhQE0G1Dpdmz
C+ZJJM7mW2kgL+Qg74Nqpeo0DeQzYTI1qxH71T3fHcs9JGY9fL3TNYtsZqofXwJw47c80RQBLmxT
HoJ+74tkHcmOmU7XhEHrXTw9+HOQjck7WmX9BAfMkJxLmA6s5bcVYztMWar0lwXR14A04G4k2dP7
6z+aYA7BF/YN+lzhCjqSFp8jnXJId2USojqW+V1nDFvnHpQ5lSsy9FXDU7tQDdevWZTniyULyBjh
v49Q5moeWeJ+zvN10p3DTDhwE24QKlHN4zx2ZAS+ZBIA5xfauQSBNXKu/orHuTgqa28nnWBGpCXh
eByc5GTnoynPpPdnbVW6s7KOcxeLds2rp+HnVAZJN6HB9XhxFdAgasoDlM2XkDm5tm8Yx81BtR0N
FUjXzCr5jzSz8xIm1W7uof3H0bfim33HBWw9WT0tAgH9WnwuZlAWXYMKVNwBAP1GQTfjJW+/Apzd
Y9IOLV9bUULrhpFN4sSuHrKClC93tVE5P2Ht5IYIysPgk+DIqY7DpyYaUf8hxf9uLwh92fb3llyM
/nOW7ZDqKsYjaDjW1QKBtRwsG1fg/BI1L1XNTVE/CkRl1uJhbH1Bkq77jTaRYndDpDUQo4cA/qar
uiMbWZ5cniag9A/QwgVLPLeYZbsQG+isJHnFOSsBtMA8kPpwUX9iAodsar9ktIdRRtIkJV3L5TV6
n0IDujaXuFi+GUf8x/XRi6YJ5WBeCplJRGh+aHW1GSqNF8v5s0duq7hstsjAvGhRX93OBh2xsRjX
bgbTsODNKABWHD17Kt44ZxxdLzxXkprWNjNsTGsXfePqj616/Cg+8mHgwx4eY5XIRwwk2cSkl+Ll
nBJztMuCGS+B29Oq0J0CTckL9IXnPBA53NooCrXx3Atzr89zhmZ7p3lImqKM6otFFoGV/zo4djc0
E+bcwiSIAdW8Tu2jeJFGcNBLOWibJfEb0GcDwSasslPKgaVgyQdlPHGgeQW9Dabi3HCiUFEEfRCq
Zwk/CasCH5ktyNBuIkN4Aquj9Re4RaBVX2+9ME98jWkOa78sZhP0j7UZ++/QV7jd8PXQjhJGdMH3
hFPjFMoV8Zb8d/+q0ancmyKCFTcyBkTljkqvQTpGuPlRL0oN8ZSILZ0b2GFjkd3JjpAH9MfD978h
efVjeRcAJlg/kFNB7N/Px0FT0qi27D4nfEr+drvNLNdCmiHUDUgrrMAPjomzaJT0RQOQbcE+XW84
qJOIby6GzYd2QfsfsjMOC1AW+w9QoNpa/VPjRJYaIrWTk9Dza9zkFj+bjiZOcJooPRcFsdUg+ger
UvVH5l1OVH64NLetIeFPpfFO4Wc4GlFSJcbXihpPCh3eDqzpAHPcZuM6JoDJlQKz8Lv9WSgzEphB
YqapL+WdHPn9uQcVfmkbReqYdldhY5+vvU4gUDKzHWRo85App0Iq0AGW8Nb7ErfuadDbVAZU+sRZ
rXsOHPPqZa4Druyuv+dYBkdsUEwrpO6R5fv8TKVQx535mkW0bQtAIK4tpxJw4T+dnEbOEiqF4tO5
msUTsvN/hupTCTnHj63bG8Ew1GYBzLkzL0n7hLPnWViubabg1zmIgJuNNOSTtcQPJYiK61Nr90+2
O4qmCtJuls7mTwiuxXig424ov1uvRS1k8/1Tg3tZJEaT2tlWzWDoUVOmY3e/jubamcTXJz6KnBF1
PkzwWpeIqJEBf8978Td0Cg9vYfDjv1bMwAh8B7nrZGOiHUXvHAPSjPMtEz0XjMlzu9+zE+jdjH76
mRa3BE8ZxJd0pgOz5RXSuqjJsYEwc6/9CPhfPcklLIgvB2eavThLlP+DjxwkVg6RVt/Y/+92sZE6
etg/atcnFeeIE/1ieDV76ZQQ7n6UJCsM47p/WYjMbZnXpAWzHBF0N3Sv4f+t1RQf1XZd/eGshHcI
cQhRmWiukkRYxNqd+Cl33oxov5hY31WhJmCqIjf4L1t/1z9/TMDzBG3nScMa7ccZS6eFxkE3itoX
zzkuGhorQxfYNmN4NgTk8WlnNBKwjP6o4tUOlgPu+pCvtGvcBX+giu6MUjDmPZmiLDm8+E3pak+L
jznGyrJnFr7SzDm99LJ+62yLAS4NYn15ALvoDsBGTYt8/IeMPrnzEB2wAs0K6CVYeVlxI8OVrmYL
RSxDLNG//TTK8KzdFhSsfYHixw6tBrD3zHEgogLphvIMzdsSwTDqCM9nBV1CLhLMRGMFWBt7lrQg
us+IF212EqzB8NluMd7n5TW+QWiZg+N5bMIQGwUJRIymBI7AO5HusUznFlOsaVWrXmB7QF94SY7N
Zec67Em12vr+JIUrZ5MGoekLsD2m1lNDFnEGRTqDwYx0L6V7tNDTFbLo2Rd7AxMM8jZ97bEirOTe
taFtdL1pJmuy8knEmqegqeo7xic+iMHF1sQCnDXO2dJF4Aw7cKWmKvU4VYasF97ABwp4sC47gF8B
Qse0T9njh8cbNCoB0TaorC4OA6OEb0c7tARY3mOWgTVd53LPjiol03w/SonwjlzBbzAxazT7Vtzr
641YictEKcJncAvCwNjRMd6CCieDTR9FjOlIOJYgAcMCGNwHK0hZVzNx9vY8wJnfEnd7fZzWXDAO
xvDqa/c74xwX6NOfZctBCQDwae4j71M5/K3+fCMwBl41UOgMsoGu0oKTzISNNLyMfU2RuazUdi33
6/f37QvpWRdkuYcPX6UdhIE6UhsRn9K7cNH7oYgHfQeYqeyr7FYGhJYogRsatro+ZZGKciCNzI81
kon+dxYu8ttExKQUFgdP5krjSnytjQ0ps1vJLVKw72v0zDmbgNqAS2J7F53sNEsiheTYuSSTmNwh
MV0tyAKm2smFYF80pT4dtL3qQHb0v1fu2KxLzVb7XYq0A20FOxC+BhK02ibCpT+Fy7GaK1pJ202h
mNzGxKyb0fwzb3ehUFU4B257quuUuIdaFRq9eRs48SSeLKFV+blXnzP/KZY+Ysquov4Z69Y1Hisb
oc0foxI26BJh0I0CnuGEaw9BK4WJ/de6Zrh44PWrn2OIUceD7nkmYQYT9nI6UYF8dE3RQ5s90y09
0dvsOwDbsugPBRdPHXY2VaICIxp0QHq2UERC+coGQplG2zELqsUN9JbsJtoWhGkbHfIRzuWvVHiH
2cg0R3TxY+iR6LG+PVFtoLteFJSFuEwTNGVigXThWT8PYv1ShamqUvapD4dnIfSHUqAXHL54cojP
g57+ROj7nGueN2f3ULl4t9zDQb8DymlgiLpF8cRqEs8GgeU9vjkbTDALXlUL7tjvJFyCGJm6BGax
Lzvn6fGenthbjyCSsAIurkkjpivTYEG+vYXuDkNsur12keBG2STViUFAfdERAsLVRZ7elrlGLY57
AYaFIPL6CHmBQnrB9LYOgZwpmKmERFW/RDGVAA1U8mrq0yZMPWLHNldoRMg+p23QlQrnNU1C5B0c
nRbEgB/ExIptj/MoVBI4FU+tiIRfDM2ZwqZOEDbTqZbB5oPMLb9eOemBGnQ1Bi8vpN+zmaVGRqFQ
4e/IFKSzZkT/YEiv/yfQBs+BEyGWrYf6g+sHnAvNVyCQktl51kc88MSIyAZP0ruYvFVXM36PrJo7
XG89qIAPDTCMdVw2Ft3otrW3IawxgMoBYZsLDhfg3eKxKHKepMGHntxZ0CsEikO0yr85hX+yPVAH
znQuaMN96bGm4H3sOzmQZ4+NPerVhpuGXE4gLqZhDekBkUKosPjytytjVMPn2H6VaOtX6jgLtIPX
UzNi8zPJao2Sb7xojwDWPcY7vpoonQ0hKV4pdMOXoCzCq5FrK5zqeR60zqtSDyVPyThbWeKgG3+i
/bz2Ymx32l0j2zGVl2z67j9PJeTRBotjlhOHmwGQz1IUfNzfh6RmZGEfpp6benXSl4nWPMNig43J
/H6Xbd/cmSeDXCVJVzowzY2ESsm91QoPWjT9TF5sfGC8p8Gl3Z76QfYJwQ4DbA5SBVPdyjjdOIwG
zrBt5svl1kkZFsJaEwWU3Fj1uKKydOpcTuZqSQxs9W3o8NkIRra1D9uNDesdJ6WttlarX78DpP2X
L7X+tpJ5tvkOlxvDH/Yo56RhFHeFKihBGwUya1YEPgZzI61w7mm4XBe7nn/rbEw7OMRo3e3ZtDKU
mXxM0YLQhB46IfpFoFTtSgI/s7AryNHXJg5g+LjeU8+bpztFe0Dj1r0Dd7VibMlyKTpjdRQ9jcWN
M3AK3kd+lHIXC0UEhAAFbjQKHTjQ29sh6EZdvki1tuBOcvcCRE9iiebTOZOYtHePL7auaaoHZ6tk
oQQgjxYu+iNGxGaGW67Ntd95yTHe6YvrzdVtzrI3oxPD/bA+lgoENOGkX4FI6YBtZoGwZEwyN3t3
VVzTQzUn5SnUvozhEzYtQ614Bd2YXd8fclKNf+m/FpkMXaOPe9Vr/o95+r0eYfG2FudyHL1p6wNP
pxSlTaDx4U8JboQeLN7bwbe6UgPjEyo2zLxkf6ReVRnVzvCqON6/TgW9j23bHkR55wA5Ui2fnPUU
UxNe/MD8WVeuFeOBIxqBfNy3XGbbw39rNhMVhJERkubJ9sxA7WXefexJmgWWD4IjYHUaGJI/mRig
6SvtINcg+aCXMCG+PSPvLLe2br2aSAwZzKLtgnLcmx7DpIc/q8I6a7fXSu19GefSh2QivQQZrhDw
5gzXOzhCgU9pl9TT98i/XXoVx0f0NByvTQ3jIxb7aqf5MJ2Jmry2NTo+Xe7GGS1FGGZyut+zjS5N
m1+uYhYsB+Q21jpmomzrF+bAhSQI3f4xbfO8OzI68LNs3uTioBSzN3HO6HETI6vOUuQUn8R4BS30
JBWqRWDZVpLEHASVtAeFmJDDL22A3rSVKlZ1zlGMOBomyg2cEGONTbnRRiqtwKXFdzJSrRpok4Sa
JrWGY/s06CO414O8ef0mzj99iEYLpK7KZh0uefGwoXaD61ExOszRtB3wVK+PJZ+bgv/K9g9K/KQm
mm32+c7MADylB0LeRR6Z+WQn1WF3MnOQFYHp8UPavV6+Xc8NdqCEm3m+fclFW4+7fC0uX4YdOWNI
OIH39WUf4H9Thl+HZ95uVF+V4XxxFJHLfEWUzm3dAQDuljLPuV3hrBiux5XQBwDTPOS0LU9qglit
fp+tFvOKGiXwNSJzZ3tFbsjzEkyiTTULRy902g7V5Yo1yTU6U6lLMp6rDNireg/EF8I7w3Z8n+hS
w3c+GSfRDURTHRslinSo1Idnkav96jHHm1UOW/06MZr3AiS/42zVb2K7KHwsjIEX+KAG8F8lJ1OX
+7X8uzN+UUIB8a9oSChO9VzRlmVfJGawGe5iIrDIc2Js7lDdSdJDfDSPnMvDvxC70+8aCnfShTbq
nKQ5xZ69rcspINZcUIKKrvc4UAS+loqfEx+kuIL3j6BUrU6IgHGbSora53nZWzCDUzDgE5Azubcf
URRsFK0/o81ZTvbuGefBeh7lJnIH+a4qc0KbM6ZJ844iZommT6/xl+NNVQ7b82r0NQXCdt+yf7b1
I/KAEve2vc/aTpUrSmVVrmrDsn//wvNC9W+ujog3UKZnHF80yGMiwJM+3adY+U6MMldQ1b1ZZOLj
lvYDScaBevIs8OdAY7MkkRJdjxlUmTRFKVgc37EWF7vUNzwJ4o7PhVUvQTRdtRFNfDgM4OoAkDVN
LjYLcMR9ht2Wg+jhGsR/CH1xKMcNHbqbt9qxXoOMdzDQTVTnmBlSw1F1IGItFnLI/ZhDQSwgC5eX
nYf/IBwigIrQHtrsOy+llZyIuNkP0FAYFJ8WJ3qXCh25mzLxZYGqLpKCv24oLrG+HTw+dUFRuc80
doeUmr524HUMBkq1SAvAVDYqTF3bqVhg2nxf5aCzhjugBHPzMkhyNMxCbz3gENu2HIJ7oyCLJbzm
PAw2rmQgRrFfpmKB499qndTJG0wXPNbhQDoAImW5B+WtY6fqGvR97eCZtr9SRAT1gJkdlaACyOwO
8HSJSFtEikcQtiAq0C4d/S3/IdTcAFmQvfK+guChTMOPkaMV0u1pNWv+d87gluia7+Q43jB+deRP
NRb4YoE7HP5TZKgJQQGi2YHBpG4Id6EFl6kjydhQetF2hNZrXiiUSPTkQJ6yV0XWjemJrBrq1b3l
w5RlgVHzGlBfo4jziyTweuGfKVIzb1OfPE+iPlQOMU+hulDpEHUQOTBnuNT5XrE2yg+RbKqtIA34
2jXCq9tx1AF4NmobICbIJwh99c96gx/R33tlmpXJ+79q6fXuGbe9sFsIRDGcPKhv1u7onOeD/NVu
QiR4WP62TdOZ8pbUYGW6QJ8d61eLySCdHe5DA70uOSNb+46JVf3zTCDOlzgrJr0jYwnyQSLtu+q4
ZLzHnrWah3VScMf78+csCCzx+Tau4Lj7AJEmnPSclqk+EsmLsY21anNXRh4EA0FNs3oAPrxmPTER
pBv+mKEEBFekLLTs/+Jsm5LqqlgL/jNca3FdqDk+DdfsSLWqYkSzZ4SpC8GQid4XyqSoAYrVoaB5
fcbwy/wIi9/HwvWV+YtB29mRNb4ZoZYwVYcxe8oTMe5Yk5sJnmJBJ006fsbcuLgfuKAJ3Xf/M2S4
XVoA/hY2WmKka5jVhPFYOGLL8NUH13IEI2E/XIjpcRCE4oPE5ERbXMwA42yQ5gGdbIX3Mzcdh0Sw
QfdxwoYudvZOYTfl5Hu0KLUeC6gJeUSovnWWCYtXBef+OrO8bVAYzEDUW1rCx3zfjRjXdU7Gr+hE
G+bPbGeCrwFQaSVsPwR+ETJ4r10wO/eUUd9vV/JzMxNzcb8uhXtXb3TEI2CORsiYwW689EnoAl2/
jZBVh5cf1phWe40bHorfWXJab1FLEXxA0SBLNjm35GKLsl3zGT0cdh8AlI2uTdpvOeYWWSGm54ZQ
sqm6tk3RlI+jD7jnpU2j5IJClfgLPaSpSPRzD9nH28eUzL9ITIduk84kVYKvJLYcFefD0tAZtg/1
xL1jtCsbX5j7g4kCqq72ZqT7rTBqzXt6qCvRqkXZVXbCnP4w6vxLBPa5QlccMgy3ex0COWGX8bSX
uj5GwXqgpihsF3Ekv8nv/wT6g3eYxk3rdqpruC+fmfQ7+NwMSBdg+TTFi3pRPYCzXBrM8AuTLZCm
+PelafQA5ZyG7YKLlMONTexGhvFx9rYTJIsnOyI1l0dDb1YN7eQMrR0qKbe39feUHs8IheWtV0nC
da8B1mm3LgqGstM5trCI1DcHzdB9GykTcg7AgqBxmI2Uh8qaSY/AKUWkJ2wCQMzFf25JQDu2ubwW
lEbX9dO/ILbCvznOKJ8GrgxvLIC404vU0UC8TAmy3U0Kn86FDvELuPbdwDixrgArEgUH1pn/chmh
MvZoBIgIT2CupswNIRTRVgAHEwd5cPXumvsNm7rZYui7jdOlffYSoAc4yfMGrtIg7+cwA2wjLjRD
5E1clF0jJpPgZ5ndbuXjUB51I67nhMx9J9ZyWPlYfjCnH1hP8ydmHEw5XEfCb53zLP/U0ZuIwxw0
Kbx/zKndXV3XDS+k/6Bba2Xl5B2XBF6/rdyazADMT80S2MVnXuOMs+X7CK+v65/JwtSk+b0ysdpv
RudV/jODtAAyGp3XMUmvMKbuc5Fc8T+lb9wIKggXpzl6udS+FNINqWFFaNPDFE0oPBCZokO11ifg
IzGAwNJHhl33N9kjPhtNxwqO51A24HVPHS2YKn7GeDYeutxv3GTxkNfu4IgTXycqIVkHkQkXbpD/
w8696h2bm6ocIJjTDstJgJ7ul/iyN3z/VTD6YeDFzHjpA71+05umSOqRdKyeHwFf7mK+sa5nKVMt
CcFz3+jP+2TSFUJAvztrQePTzg7C0ofQMG9JMCSDRxcMiOX3tP4lAiMTgN526q4d4ViY7GU9k5/W
KwqQQ0UZVM2zB2FqAZS8Y8o6Qiuf3aXaY9NTNmRQp6aNTjYZuIocVPt9iOYWzedXATVVdrIfj6fn
CLfK3pAJcmneKOHuEm8mQhH1sPSj2HN0ZX7RmVInYOCkpk0mOcYXvxGu1zAWJHO/mh/xd5xU3kvt
wZYg/q9cAmCIibuPuScctdwZ3bDjAd5O6zGoXy+kCfxrDSyhnP93Es2W7PciWE8zWoUV4i1X808Y
SL+N0GGao8TvJzu4pfCDjsQNdKCQwlImofPjreoZBw15/hNiDD715dfRwlQdGiajAWooNeoZpOhW
LeKcORrm6wilYu/1p4wvVNUd7oG1aZwMnuXguWSNTDqI2svM8h8V/E1FmmsA0ScC7yzLCcQuCCQs
KeCVMZ5yqIEuAEc53ZwFfBmrKl7h01pvF8akwBvN8rF3V1gPboTVeEYdjfLNlXfmIgX7Ctt5nhVM
FHbN60Ksu6fkO5lsBhDvkbnUIXyL1Y3rQ9BJEsg4snIJ7oqNYgmfxEzRuempWCPdwdEEx/sb1vSy
mXZmLMqerFvi2dQBYYnuWFduSO4x22JepkuJHfPUyzKuNGLKu6wrTZt40n/DgNROSLvXnA7uN0wr
tsowf2h+e5mYr8u7HF6JrmH9y+nNjVY4wnHKsqT4CR2fEgnRxXoAsQ73MzmpFT+QFfqWo1XLB+pg
Kj2fx+0pHREaqnwkH9tHmvvHhRVXIU+KM4vdHsr6J4t5/OP1OC4Q3rWXFapFp00smllpKd/ClMRE
ulf8CPs2f30McQuQT28TDJ/RHiWzpt2KQhtw6gqdaHP7VwIVf84hl3a1oBPHz8WLVV/STgpdbyzE
0Qv9TcjugWkAsibMSFzzTozVbn7MifRXUKeD47vqjEV0crm0mROpPNwWiLwpg5/hiu2j3e15GOBH
nGavVItOGSguIxXVciRLSRKU2l0TFJxvUPFYoq+auvFBhvzxBU4L5DTzuONdwFaBKoYKPeJudkhP
kgPCAlZ/n1EzX49qXX+PrBulK0VeVW8b8K7KCuSsv6CLpXwjpe9HBfYFKLcGb8lxzh2sJgtRCHgD
jxaqHSZD3I4AY8fRs63REXyyxwXXPTp/DM02pCc+HO9+3kc2huooUCyXi2B7XjS6DhIZY4cy7RLT
ahgPXVnY+Eo5rTXx0xoQfEKKaM0wap8T0aE3bpvGaPE9z9tCrOzM3m98Dq62rZCq6A2PGuazIPLf
qpbHZ6synjOvECvdE2xFf1dJMDHguiNlMZVFH61c+NMFH+Z0D/MVyVm7DNXqQavpiTLra9XA9PBp
S0D0CLpZIZBzsn0G0wo30LuT3UIPrmNuVa+jlSPLR0cygjIYTbPBoCwveURS7vP6shcrNYzRTFWU
uhBnCeydV0nmvxtJxRk7tybmD3TZSMJ+MOaLM3wFrzoq6fnX1ztVROGVKBGAx25D+jSGi9rd0VgR
C5bS1FNByzLg0KNDxLMaxfvtRO1SfW+j3c0h+jNWNA+V/JqXwdI2mvgLbNvqfMd8wO+KQqwSUFw0
IJ/xwk77zOe3vjOy4rVVEpXpBoXlbhlkjZpOJD0//mNGDOWzvg2R6B7++Sk68Zz7yG215zqWEp2V
lv1j/zF8db8FCXxEgdHBPFZ7XJym6Dtfn+2N6yxRVbHP5uZufPAjTTneJdXqyVW4K0pO9KHI1s7T
AWQz0F8fq/jjSbXgeZSgWQ4ciVWDWTi8JF6dSm7rM8U2mjfDNckOdaWqa8y1nqPKmWpaABVnaqxw
r/yklP8roPNKzjnDW+xje/HQOs+RilgfkYCpoiA1qb7ftMSQF4MrlPo0SrnmZBDwpnjROwqG1Tt7
hHTyDgc3hx91h+8Gh3NZzqminreMCPb0FnGy19jmGFlsz9/solfy7WVptV4nmxOtWXMQsNzXexdH
Iqy60rjUcAUvtbeqWYtirm1oREKWULh8PkMZ7eO4mpnL7FXEqn16nX6QDPpm97YuQ5Itg7vgE5nQ
JgPS0oGiCZvd/rylhDP1ioVWnagbpqt1ICIPXXCxrv/0wiYEljCFi6D87YnNHa1ffm5gpPBlgqUL
68RqLixNUFhvH1oU2CA7vTX/Gwoab/DGLWW3dDJYmAdSNpILFAMZEJFRTzuTofluJHb08XIOhyF/
fUZyiBzoWoDNZOuNwujNQ6ddA0lNCqs5NYeqO7ZR2ixapjg0tfQy6BBHakXc/QiT08V5YValQ5bG
f3xZgnEkUfbgGQn24Jl3IpW7kr22NswHEnX/O7533xlPrvlUeVcRRDLyHuH51H7a/xUMQtCEivHA
Z71qVHlukf9MVeSfHLrw7eytRTmtkRozbCv9qanpqsaLGkWtxr+21bZBn74yIEHK/GBojusWjjtG
iO23auBgAYuTAyaZfAPIai2clYuy55kOJja8JjOycrq4+pkIe1yz3RpdY5yPUxPFA03VHi5OqAot
IZhEla/qSERiWzyhmfhHXGksnkYOImfLg5jcFYRAOdGwMtckVWGdtDjb5OZqZNteM/3rucYvcZZY
+GZrcuTvhpWpuUurCKGM/KtlIxGfZPE3Zv/rACO3s1kGnLfEkZPkCoyFWsUC15qfCOjqFlNQnwe2
BygsmMOKPKuIzi++OxAlzATDLocfwndS+EzcAxSJEOHL0xsphMcGm1yn0tsWMTXYkdtD5DMAghrl
BiW0JP1IoaCT7uHSnZwN2Xs2ecg6O8z4D69Y14/GkBn4iZLccYUd+qXhn56UAoSl0S4eUmVa0dZ0
FKTPuzBHJFRPwxEvp8K1DCV2bkneGcIZcH0Lu6fZ0HOzp8hGGF8LEozkNaP/trKuRgq0yxU/Z43Z
KcLxmoMHdBhxXMoT8KAaczAYSSsPCazlWwiGiBz6UKZytd6BvLssxo9vbt9AzG7//JcouDMA0sCg
Uz4KMnqumKElRoDkJzFjp2tMaPERpimpxFiIJrnO/8bO3l8rTxiUo0FGtMIh7/QgxmdyJY/M7QRZ
Kn9GHy3l0ZpY7zVuYtHjC5gSi0vpr+je4LnZTdURnCgQQW/lJTjebGLGYrDaoy6lxeONkmGAjpSc
qHKNSGRfuECKdc+pXmEXNQ4xWXgGEK2Nzg6dSvuRr+5ePQ8s27Xsm4P43EfgVLrYwK/ihIgil9XO
3nmrUnLZY5zGTtowTPj3BQWiSTLcdorxcGRTBgQLnX6TgJGDMd9TlM4OdZmorNtUABgV9Dm2s1DW
/72WTdLF9qom25IqvGvmkaq2P2hMCktQUqXB2AuXevi/xwykRaamWPY/uwc/h8BzNy68v4x6a9GH
Ad69wqKruTVDHGRytLH3ASAvaCJ5pzKV6TJKVEeoEEyJe5ndh2GtJnXURw59wSLiaPF/i8c/g/B1
OtMMwWte6PVDZLkiLLHGd5/cpxSmCVq9vlkZkNUm05RZkvMHPrtNT4sUyLRf9gv/lXoBFvmewsPP
x20bYyjTa5J0aeFQT7T3Vt25sS9hfV1Ea594zZzFS7ejybBzOxpOXmNZoIe0aMhDqiyq68HfPx8O
b6xJu8UxaNpsmB+zMyxnlo+GD2vB9mVMU9Lh3GYKm22xw1aVLHNv/O0NnpaibHv69EXLpEk8saT+
4sXYRxkQtXMg2yICEH8r9vXeHGpzvUtT3TH9X8dlA7qrBzI1Qd/7WOO1EsAtjLBHWfGkv+r/BrCX
Pxvm6+vANiavBUIvIB81L3D9F6SE+gefpp3MuzL+alYyEuC2fwPBSvJPtgGAhGvqToMbGE6B7mc9
jvhBJsaM8WEQHhg+CYB90E/TRPGQ+A/yqTJavgBt8X4OUgwg+G0Ix6ITp6tPQdyTUFj3ASMmLzYu
sxQ2bMUtr4NZvtenLbH+SYsvMkfrA3NUeHEVlBtIMyZFB9LjGXPYRUgpCc9WCR8XdMSm0lPf4zbE
IrT/50vULp8edBzNt6XupJkkeELrUiLb//XEpncrCIG7RBmhIvNjjk2pTzoLYL14WPzgKqYh8LNO
Hup2RnV0ZUuymdu+VDYwvNwUCsVcNftYe4Er4UN5YEN9zYyM/94u9WGPvKdDDtJnAqtvyVMy7RVp
XzxFx+rRs9eQoeX1eLMqW4T5uew4bgVCzKUK6JYlh4WxSEU1j1Gx7Dz2+yXnPramOkmOfKPQNbEW
/37oobtYzncLhf5YY/Xa89Wa6Svj3b33OTlYb1wZp4Q6poIzjuCEMI2zmNJo5FokC5mzoxHe4Sqi
J+EmQo3B9HXG/YlHn9gOsRj6lN4gM/F0FqXtPv6KZWMRw/NBJRdp5YcBB1dsxfGXxBPge9slikq0
ixR0SLPKZvTnSULKj82hAMeEjrUoUVCK4W8IDuKYP7U9+OVF8zeJ+zGVAVInuuiyqnPvJobjYaUm
Cvn+G01rk9F5Z7c1YQvlSSPERJfSaYgZ5ibsdDlYMcxKQX8z/1dMEyoum4/zp09DqEHFw2ZulcfR
b0dbdd+NXT2AKIK79folqBkbjagr3f0PxJlczTxJccZ8rI32AvzJn5ydn074FF11JqmFtf3BClBg
TkJja0XyNHyN6/BhSSoFYQDbNjakDv94ArspllZAAd30gdP4Y8EkI3S9U8Hqftiv0UMwejfpWCOA
+QC9J5aAPSF+pRVympPI1PjmE1Q/RGAtcsVHAbB8FwyKH2u0wDQ+rwFeNYVVeTfEZ2omnpXOSDzf
WU4OGJfFTzymrSVzBG7bHCAUnpp/3xW+XRy91vldu6j5672db2yMPJWvaVgE6xWjtpDF8b7og55J
apdU8Z7vlsHXUcqwkHIjQGS78oWCNOltDoAxQnJ/KLctrv2x59OgEI8GcQoSg/ImDPnZUf8BaL/g
un+M4kU1PMSy3eqshQL/SeK5iOOoUpOOvsYGkklYfMAzg/GcJ+M+UsybeyaAZwgGjx06vHhZCnPC
NfcqV5HELtaXSRfROquXsv23trYHq3x5TSAZeLjojlpNA5lVNGdoeJrWE4NtNCQReziUBVkZIP6j
1mcRUqFVzL0MsKfOk9Nm7cp/U3EqwaCiD20vYvMznSsSW/OCXg765tAV4tuUnysj7QMSDYkLi5Et
04tp8QNLn5n7rCOBAczTpvmwcj55BONX6xK4eZG0a/6oCM0cCtKHRlQBrsLA1zYbHG6Z7CsljbwR
0EHfxvjNyLn3TsJhYvgpuIadiKxJvYYRZ19x+51xkWgeKZjRMT/Ei8sMJUOa8RtSEpDZC6Mm+x2m
zhucCam40vs+zkV6lHD5TieLSCdJWWPCjdg4qok+sasSML7DN+Dc63qvNc9QI6xniCh+Isk8oO+c
KJJHEwEIPmxegMMFLoqiCJmVmwNyZPcJXo7G+HI9myX0b6oyq0u81dlVKGeauqVlGixfNBipYik1
g2DBpbt0fd1jNgm8SwUtHhoiN8CByagevogAVfP1fCSRbaU5ukYOr/KKRf5DjMF0OKx0y25T+6yr
CnmHMSMFpJjDUBRX5kHp2YfwYUAsDG1RhjGWopM+JUALxxpFheS/7JvK/L9+Fkq4jnMXfikkNVHn
ByjF3fNgoJIBNExl9YnbY8Qb7IZNBtOa+gZyqLd4mci5YH/eCsUl+v1qdv+HguMaQUc+zUh4QjAS
UoYJQk/78NvUFWCnRyVxO4q1YAIREdWLF288BGL83wqnirntU0yhWnTTCSKmC12acO1GdzAbXueG
fbsKO41Ori8AwppTQtbkqjgddXJ/DVdKdNWh9alsLKXmtQUFIivGCX7f9ajLAGSaGOASG+SIr90x
s4wtIXx7etNwjZtzppk+hzXH9uQ8Bal3oF3TM2f9VuHSG3XFgD4GEo7fTyqI6D0iWCQbtlY9Q+px
cVP8tzcZu1k1jX4jpSUXw8y2yVGAPfye/qW0SWGz8eHa870J3lGBShepGNXj4t2jtWiIibVpNC6S
32zJ9v7jGK9SpeCJEAkWkwj7DCFEa4GrYt/iFPhJfkTtjh9JLYJEjNmeelaql2mYLgQ9hxMxMUX3
I+HWYxkUJT34rR3RwWAaWKZJsfhysoXrfzHjgGiHkqxU1d4KL8ZG56FLYr3e5qOr5D/CCSiaq8CI
bB/5Wi7ZHkB2i/iPWYYQqUt3ydHO+sI6JiDK/FZxAxgmouN3HeZqgdjlbM9Svs1+Y0whQTU4XJJw
OtIsoPmzvYnIbCCN0ckwtYNzVCI2kNjhAn5ILurzINidOZ8EwEkNLA2avDwT36eXuO/Le8z9qau5
KzLDugJPBT7NFOfvhCIS4aRW0+BETe0p7nlFa4py/9rAINcChmUc/dhwL5G0oXnVkvD9uFEYasv2
VqlfeR1qIOjzz36I0pp7yf4BTq1zlVxGsW9LZHnrX/FAfPXnxlMaL12v66U2dRW2XzY3eHudEHfC
dfePAW9KGXi9rhLBIHqemCZD8aiIZVN+Gk0phRkpliQkIdEXH9GC5WWDUDMoigoteNDvEVeHIKlQ
daKqfPTkLEKQUu4T+hJPdlRg/isMc6uV34DwgLFdR1lEP+Zc70yr+DjM53aTX8mEvq//JC3dlBgh
n+7ItdHfR+0XiY6dCjM/qFxz9FQcHJPiisy7GqSGgTM20HhE86ZuTRKVEZbNYvZrY6/P0x7iypGB
f8/m2E5Na+A8VGDmB8lmdZfe0i3JCSSeP9BcNiuYAY+byf+LldpQqhxcXHdLVo/0IvHtpRdMNK7j
5BWKZov6+i46L68EYAf9ZcFVhwhNnt63JXAC/oWyyBvHUYSDThNRkTQ+P2KQm91V6i2G5QepFx+S
8at3wfzmmYrX5EerVp6yy1B42Devt9rwoKZgR6r+moMlvPnghlQHYsPtFG+zXNhfc/MPQxER8obd
5D8x1dFYeNleVot7J4Easc6sUxcqr/wCG6Tpfal3q5sGQ5KlwfWaQNi4ooawzck3BhcWjyWzrsO3
oHeqHAbF0e5fIlU9QJEj0V9DcWjWxCv1E5B/oWgJW+E17iWm/ijLTLc+duKukJx3nS7HMJBRi94b
Li8nwEkAA1O7azczu9H1xdicrazKc0cacyKaHYzSufIOP7JkzAPsv8VmuYQuPxNca2cO/4OslPvt
6j67F6qxp+GzcBF8VRcxHMH8M4+QshHBpPfEj75sDf35OwxaSTKlt+hIL444GOQAb05sske/dgg1
3Nwh7NYapRWBNhZlrDReaOaQrX7NdDUVnI/OEkFyB6J8Pn2Vt/RbDKFWo2OKK0JKJcGBQhOva+6e
omaKmcCmWx8130tARj+isk+PyH40tE1BrLd62WnAVw4MhrBiVH3PC4rID9CXajVnGE6iV9wCFVl7
MDZX61h99bsfyfKIbzRFtURM+wJNUDppzNMh3+9bNtNce58+GvthT2QF5fSWw1zQMG5VtF/YmBdm
7qujHolS5mOmgXLTm9U0oj66HjnglO13h4H3RRpWm/8JvLMYD3fyJFrtI9YP75Q/F4CC5pL9kgI4
E2HzvKrcoVD8erZSiSkHdA/1FsC7ly3iDPFwS8mfik0K7L1lUtlA2US4NX7ShPWXA5vTPdJ3XBQ6
8yyRoF587XIL5IetjSLPVtePWZetFslBXXwA6+7Y0FPp8xn+DY0RbC0q1SBdMN9K0VKZMZGKkE6r
wrYoD6piKAnUgblCHjt+PF9gBSRKb+v45NCsj6zhQ8554EQyLQ4i8FJlE+8YyrQo93RW5dOqhHNV
91euFvIgryPwRSkt1E302n6rOTIfL2eKU0Fg4/i3AkJum8JwRoPrXz/PCjlm+8gwvdxAVk6ys8VW
Rv6xQ18P3wfq2jX6DNQ4mHyRtLAYNIqTCYu4vgWi31CUzSUlELaR2kkho/IV2l6eTmpP9t/+jNKc
SjGpXxLOFjWO4VMyjj9+77jGsrklkjl3He14QG+udKrBrPMN456C9N22XMwJwNbrfEY/nmgthfnQ
uCzKC2/8k9cHm3uOVzKbjKANyXfXdgMucUsz6cRLTdjq86gTNXN3uyGirz9XA8iwwuAo0FQDOEAI
ZTQSsMDOWzzu+EhHdEU7uyPuuGEj2Eq1Qb3LgTuAqrrabFKMIUhD+Qmn9Be7b1AiKXUnBi4wykU5
M65BGY2dEe9ZW5Q7L39+84HKw8jqm+EsoGP7Y3eh29MmCSsRRsDG/boPJ9yd/Z5aMgkbXk21m15E
qnusDzwGC182NCnpdk1ldBA9uVjL6Fip+O1HmnmGNeGQHuYtcNBJTO3BdUpYQ5jfDfF0PfGSuwXi
MxIs4EcorwjjLKPyfSiuNpOh8V7jTBswcTDDlB4dbWjmXXhPEboztwI9uhlPbawlYPSu5ZLzsR/1
fuiJV38qdV1H3RrtNHiupSEAtGXSaEBMHjG/bliCqRe5RDBt9tGS7rgKq1NXmQo7qpG67U/4N9L4
fW9ReyLDO5pNl2ST3M/1pXOHa6K2cWbjF838gd3W09QLh6TRO4yBogWok+zMdBbbxJIU6u1825I8
LPwY9wAPkYO73EzZxVlcz/ag4eZ09EvAffvHYGsF4tPwgthXsOO6nMN6yowJvXZrEA0MWAFJer+n
dzm5VUQp9W4VuLekSLkdGlW3LkxdDrwWDCUvRwZqwzxbj2ljIiB0eH02XtTaHrWqNJp4hzWnxB2Z
1Uy0voSB26fW31NAhoE6cLxi43ifSbtFy1PRoPVhwQrwOKqMvcfFLBMeMK1dYVg93ZiUnLfZmkVv
54hKlP9icLUqnTsKxwfZUNOZz0t/OeT5VaFJmsGyeldEPCqWhlMUZD4sskGGuiiwVahrwltGwu6m
eHf+TeSWv20KYPLIanTtjrXHs3QokaixA2RCD4rYs5cCQuOTvaygEDjcGEgpln/xwiVcxyGtr32m
wSWVDTwK9n84pO8UrsOra4y3hEzuVh9U3jO93m7s0ZASU6LvcOHQdOz3dln6k7liZex1z58dag6N
RyK49pVEkik1jMMfAg3E5uzrKK8V/0vjjLaJyOBQ4M/BWwdn+jy4pEQL8NZZfQodUNaC8bcHdUvK
49euFd+FbVf3UhmY0glvv0fsbsANFxMosmzxiUUSGmdZay6fSIpKAQ6+DQ/mXk5yZLcxBitUaZCn
ntyL46wMT/uwOF283VJfI0YIfSCEc8sxH16pwynBMVrtApfW5c9Rs6cELJfQGDnmMWElpa8T2GD4
z748ALfR3FsyTCDQ7fXdE3BsfowscsKvzYZmHLQ9oirZput098ASZSSJXDtVhDvk2lOizGIYTXS6
KclpzIa9MaaV7FEPEQordygolBHCXNDBmi+P631296gulsOkEUxQianRVndrif+jnELgDCeb2l/R
J4ujY5s8J4iENI44EXxedZKyL54TWY1FHKvTORlwaYpFZ/UAZn0sV3cijya+QfsJSjiLVicMCWqB
dBgzZ3ImesYUgQ4p1EFw/ZGOXMGTMSx75HP9UOOnGP/4elD2UCvdsQbPT9NOa805U0BmHOIyTki0
kpf0locXCDiq2rK96I8UrhT7ERWdNWLT0TKlV2j+ibUGt/++Jg/szcCL60cB3Py2ApVRy7FJA5Je
c2cMutv2BHHlD1oRH+V09O+wdn1H+i3AFasvJYNUgP1DIt+wKGSnEC+ay7/YX2pmHyZ9TF9Xp6Wr
ZAr/QmAmgIvsHh2r54QZGBSdiL2CGzCUum34SdJd54EHJLrh5f8etuYA8IaSw3Dw3ez1dYgwdWuS
c1GgvBSevVcw4a4AYHZ3ymcBedXNcOujXiLJd0BS6aUJB0iE4m9VDyzvAieaI/Ziwg4WP/Jw5kuR
oW2JbylwHRl0C7sVq4ofHSljYs6ByCo2PfLuOam7M6p2wKG4d0lLRP25xf653jifdhYDluOl/xUw
P1U5waDdyJQ1ia1yu7F+XbLBucBi0nne92oz23NgMNVydHTO7R8Lvm4qgRZ0DUK0Yey6G87GauPY
rQUoXWdbacgE44Hr7qKDB9m4a7uACAl6T22B7ve7ISJtZYcOZWTUo+pSgLfjnd7QhB4kIhb2DpCV
niA1WLcNLpytkHpndRBUlh+jWOr3UiVqukbPdJEzZoUAQyk6QQBBKhe05KXnG7UjmaqAe0JMRorH
7RSDseQ1fk0Dg7zCWSNDX9MuZTiy16BksH2mws4CiuPQVY2TxcWDC4S4YPAx8ULEPAgOrbIUJB99
867y8OZeOdRV9vE4c4dAidzSFWEnUZxMrV7LVJNAaWQgcAkxBbp5BwirSvH2965c0U+2EkrfzEIb
GZM6SSVQ4JX5koYY9xbTPVqbNxz6T7472pwpC5gG4ksLzKBF1M3Vtig0lwLAJc0DbEJ9R5SKLxj+
QERYmyYqwfJq0CcRsy4HU0HcClcHz0e5n8m4R+u4z/Kcv96Kwl2Rl2iH8U5ggNvrs1RRdETD3NwZ
C6Byz2At0qOLjk730tiTs5Vvu8WW+kjXU0Du4/8iPExjxKxKgfqeJ4ZJXgoTXc6zgdOVxOCUhZ45
LJpqzChSMBYloXEpzOa4ydGC5ya20e9SjIT4OAIxcPxpbFpGb7Ppk/Q5UBaUvZ3IqioW3rh5W3tI
HI4Gqyfh6V5oxWWns4BBoW8DUcpBdFVkHmyIMWOpZ3Gz72LiWe6ks91HPdMtciuGFWh/LIESkwGU
0sMN7mDbOR4oLQhbAo3TyS3dArMAzSjEU8wEJ8fe+8rg7ZdCSwGDFaJo7SGw74ul4VizZfHNlxOO
SaTD17a/OP3O2312eH80nwKodDRY5eeEeRmfbTXZinrT6evuk6v16b73YG+B6oDE8Uk0MrixHhcG
zyk5D2AL7HSLoOhifSDmwuA7rcH/gTPWi5rnweg2LpxkzHLcCxqSGEeJgUkThdwSOxeidO6w0ooX
Hf/KnC2cLcyaSxAV/WOkn5+Ij1LR1tesBTZTxM3+Co/35fnuDbGAGIfc8rzJj5jWNkM1GagknRCv
itd6Wuc9M1TJYcVqPf7x75EmVONfgUt5aH1vMImBZIbyWhfnCmp7fQJR2PJgBqIuXDGcmPcdX6LX
aouTKHlxk520ZhI8PIzO+mavtBgbvcUOCCXMIOkvCuSh9b1KKpGjZAh4AwnyC5voVs3IdbsmKblc
QF6Lu/j8LsXweXHlnSvBiUslgSPwQjLkSKYKOreV0ZvGZKBmmsTjM2uawFYxanSjxpg59feXQpVP
C+GJbJ4MKHLYGAd67wSHYTNjMniUPy5ZF0wCnPQK1ykNzgWBl/eE2pfPqFajrX1fMOUVVDv+jw34
9JS4tqfeOb4tFG4jTB6EAd47VWK1YuN2410qxrA0ZgnALp60z+1FyfGdAYzT0smYRskbq078TtHj
vbgOzGQ641ZsUyi1uklFNLcWTHOzXCKV5ZOe6Z9JR4MNTZTt0pt3oRnV16XXBU/j6tkVUchRA0XQ
/wLQE8p8p3xBiK5bAhvdUVRKJ8VFqgEhzQW8pJqjWg2c3UHgaAITfggBlDAPSxnUdVifJr2itRAv
v3KPBvabGrSsUEbbe8YaSiOhm/e4bUTK6aeNywcFuOqlDLFLtb0/8ZvOkTOPEb0X7WgWJukHKrJi
HZ3jWQQXqc0qEPZWoZJNRG3Q5mXl/1R95xb+RXr/s8mAhVv/Xaf7BN9HS0bfWJsEG6DhNSIr7Ouq
rRx0z/+0XVLkVGbQF+SAzs1QPwCafkGs2zOlNpXEOjkG0o+EqsGVzRv7ypjL/YKwSe5JTOvwOHJX
j7AP8dC+kFx2OBy5BSrdPOvcYjGQ2T1uCsfrfYT1PvoqTPji7Xczbhs5ltj7HRFAdFu2eLbL/phv
hyaV1STexkT3uI1eVYuHtzhakmJ+/tGur9o2rMFin2DMihBCT9WiZmn5IJ2IMk9ZgotCjgflQWEo
iKTzbcXHMBZDKvuaKEDvDli7h62T3krKwq9/wjsi48g+CWyarv1KEEOAwuc1x3FJ/8gMiix1AkzW
VIGIk9luyxQIDx5G4qvIpUltMB/4VyNqy+ryDtJS7MIhhTa0Yk6hWwiGrHWTgqQvo5clI+vLlAY7
Gj1AzQJ8UykUdzQfqleQG4Sg6UQfwHZvbm/cYBekuZqOlvUSBkdva3KXeZVukoGPfWYkFa+63AUI
kbmjD4Dtf5WwdufNZ6zNSzGRlEKoEI7puN+/GRSo4ijVqfwXKATvXaHVIlKKW79k62skPP9GiZ84
C3f1giwIND0sNFcG7VmNiFJtOk2Y4yTQsSuCKVnGyu+yqFUAUfqkUaKA5UPN4DYsxt26mBhryDBy
Z7bHcjN2la7OOYJmEa+ybTFjPsOGBmI60l9BGZASTSYNB04UwbGHoUOZyCZvI56xaMQLoMCoIveU
voSD7gtdIpp5mdDVBbHtuirBiewHJIuPmfFijY0h3CwvFlAL29qcjM1NSwzqkzCSSpV1ieRi7b5V
egGc2Ey7CL5nnyTO0/3To7MoPTjXxcem0MZwja+6+//XwkqNhkOQF+C/BZPvYLE6L+9vGT/bSKDz
blcPP35T5PR22FE1qdMZ6fntJ9NjULxbCzRShtLjDDWq6lp2+s+3x9Hvdn4WW6W/zKEYEE2JnBJz
FxzQJwpLnJACUzRT8x3IAHGcGgbtIYe9SvKg61O71jQj7Dc753icVxY9OL7gvVsVD9W3QZKisOfJ
sVdpN0ijuyevVhIgTW84Vx3NHS/IgHVbUIsnA2YoXvMa7MOGmBBkQoAINewGZ8wIKkVO333tpFxI
ytpvsGT8O9HfIDxmiuaMA1iCsCsgxUD4ZILtjfZZAc5iT7pMFmLuqD8I1EfdUNjXuDam5tx/uRsm
O/YWUfiqk1F7MNXH9yiomlDpRw6cprr8D6miKiBjcS6aIcBQgDZ/IvUny0sa3GJXNtDEZiBzJtpH
XoHp4ASaZqsBjEWFJ219OOI9dYw2suWjiUUmdKmVkqjflbL62bW4zpHHHbK2E/0hUjOHnJ5Q4+Wu
ZZ1gcLRHUJbqP0gGIzlX0GYXxCXjAF3OQIhPsLJWynEauC81UlS82EdkvRS+Y+g8dgk5TP0CtKt2
7lLTU2V8b4eqB9tDilYz2YTzFjsWJG00pnD5+vW1HxaJai+7l/w+C35Ne2pmbXe+rccvCsONmMgV
nhdwy1Y3UpK6TiLvLqKBqmQFmEaEFxlECrGPrt0Ar55wSLdSsMTGCJRxAv3F4txlwpVmUlkXkMxG
GPFMiHGy2EwsisYoQ9mRdiVUs8L1Ec1WZxiXgIsfVS0j+7h6JhkVddXKNmf6A5gUDElngD9hfXok
AyeTNfLIih6c+PtZmeTs62+1kyz37Xm4DwoI+hb85Q0Xcdd68nZDe2TEYO/FQUbaSyYnNhj1MJre
9vWn8rz5ubPXEWo4fWG/9cZm63htzIFZMhQeEZd1NLuxE1JQLaL7dtPCloJCxaJe4SAuN6/+utKR
oxZbzZ4bGGhdQF7GVJSqvY9j4a7Xeojx4KcOfveVH6bitk84qSgKdLSs1FF+AR3bJUHCi/P2fy4I
iFQZLsfn1bF9OtjoWLhz3If9znlr6mztXq2u1aFGzZeiUv0pgiQmWQqzogjW+iMW+M9tw1wCKlvQ
OrbkhFe8aBcMwolS04zL72ZXmWLBgO4YEYpHEjo89AIx5VJR7HXOpyipfzqKU7cBXGuK1H04j1l0
zxPlFzEQMBvd0SiCA9i1cdV2prlDiFtzJu5aICrvA9xjtQmgApoPeST1FBqd+T9MHZuIrEFrQXcO
wQwnSP24oKzvzhkQXufo8iliDD7bxvuqXmrss9eUHEE7iJyBHJKZ97OlvV0ErSDqKmX8Dwnu364l
rrlOw6L9FCOSZV1lDS6+qD9gmYQrXTdCtTwK/fIp2QJkmYygUJVpEPOSxBDLCgQSrUcUr5p1JMP7
0kHmIcb4OQ0SV4PX69pUttdfXswUWgBH/5x7z91rle0UtCIZJ8sWaxbKD4Jym4kbq5zbn7+VKMO6
e7gsPF2KjvVXELqC7Ug9BICuf8qxu5N9HsqO1Vp6Dxay0Inmj20Qkl0THHFK95zZ0eznmiK/NQxZ
+TQVC+ijLyf+tO71gyYjrJrbO2hlhY6gCfOdQfni/R+hXKcUuyvYSGEM80dcvEG0nybyvc0hkELS
h5Mf8hN9WO+Dy/DWOHB+KF5TX3Dvbf4etWbimQNu+1XPTgXIn12ZFlR0GSwKwHKT0oQDP6KCLUdJ
StH3D7+625AilxTTlN2zvEuIzsN+p/6tM7S/7p8wGDl+JGAI/GrkPFysOnzTxT0B1dAHtK7uGZzz
4Ui1Takya+FxdVdGeUE7rWIUuhmaSEQ36zXHqjK7tSyc6K491cHNN86ynb9EV5bmi0gx+n774wKn
Cov0SmGMkGdDfwzIfLnaO9FMespAUQqN4e1zyDeCAO4E/vk8TsSbTe/go3OLFv7t0SR7DZqr/sn/
LXE7yjtJHyGj6N8lWhCTBoMaGSKbX5FTrFZpgdkk7+wJF14ujLuC5qsAZcjcAIZi5h4BrdO5oxye
oNQO+t2wQ1crUnAUbHEbEXboqPIXal/VI9AKhb42oalDdZpZDMmuJ3bsuilgU9TxzjTmRw1Rp65q
DbYeh3v+VDv8bYQcraqNQYTwc/v0uT5O6gVzIiXjNUjMhRqcbtzzcZdMGC2OuP6yVUznTd3DxiXk
dJtAT0lckreHB8TUQ4OeDFNR4jkWTnzN5y29No26F3osqULsJe4pbcSvmYkuuPKXKsvR3hwRIOkA
YAjQtgP7piofW6xsKYJA7Z+t9MOBudeZANbyTFDRhGxw6OFretNWDrnLrrmBc8m7HybZ3SjfWOJU
Bb35Ywo1J1GLCrAxHc79ZST1r789dUmSiA9ROL9mZmEoaqRzGmD4+f14jiKjohw7D0bQnrywlepC
K+82uVA7a8noKDePfB7YfDLxqEwRfiUij+3JrKDAIbJe9c4qkcff5pfluXQG4fsrVRepFu0uvJnh
Uxyadz8i0JcaJUdCVDpJBhJoDD/IC+bmIm1nQXh+CRWHoWRBnDqMzMkR6ZFSLbUW058y1MttVKBj
nH5EtyaeKaDzEYqiy8qMabEeDODkJniIeBBJEqFOEA7elHxAqDmrTCkZgnL3slEU5KW2nbmR47iW
u66cZ8nlkeJ4TqEDlgGl+A0jb2jT/PQhkAx+f7yGyT/Lld7rhFgmxyS1jCGC5rOajFfmE3m/wYNK
0YiCW2Ip4aFApb9cyN5o3xa0JvWZpWsdBx02JHoKGNAMQeJbnTOCX5UnAaF0ZEh0AadmmL9Co3uV
6lrLjKQ2jeZ5fj1sPQSDK41CTwtSa8zpTtEuUtmpq7VV+w3Pqs48ZVwMxfYwqL6V96zWpJykUmE8
sU8z0VIaVnj6SgyKFSU4aaRm60nRhhYkN9d+7UoRA+9wwlpVKsXWTX0vu1E6ux6TZE5wpncTFZZS
CfsRrHhpVIxg5v1Ko3Ik2iX+AMZPbMV8fkcKF8Rzpnp7q6qnSycLoLGe0U8/rmenxg13g1zDvGcD
Kmyei5o8H5g2FFOR/bFZGwCowmp2Pbeuf4E6mmVAvRJNkNtitpX7Mi1wDBV08afgo/AI/kosJwFo
ZoHWCVFFCqY6KXDRirnKS5b+B3Jf/1zfGEsBv33HT/Csazn7uVXmCqLD2kSTvZFyeemO0P7iewlb
DETo5OjraaGlhV2PuzVr6lccn+s31kYXOqv4pUAYw0mZiwQB2C1s6QyWJJvGQ6NfVPWC+XcHIGrG
UIqCQyaG9ATpIk/32MjXfoRLI8cw/v5kbrBqgvUumOQ3ZuuiOGMpl1hJ2e1J4X10f33psSuU1Wbh
tO7gqhqR5cIp6R7UcxPaN/GStt+NVIBr/GkQ2cEtmXzFlmNMt4wA6tfBWhQ+iHwfVGoi03xcQK2H
hkq109EEcFdMo3M4N0CjiDLtzx+QUhXpsFm21tyi5u90BNAxSR6sIbE1L+5suSXp1B2TCMY2kijm
+DvkObidaSnjCEB0TTfuTTuIvwPaqwy2uPrRU6c8jwv+20QDCf/sMK6SSsog4yElfq5U5XrsPAB9
80wl2rQHRmCI7DFgShWxNqbMtUueTboqzAUgylLgWGqHeVchV5envK+uY4buMvwSTiyXAqm8naHV
fJK3QLR9JLiyBBl7P6awlAq3ii2L5dptP8dh/1w0EaxeH8ceqy9dnaRx/XHHhFhen2+yC2/z7J/d
uUGEX+q6F3DskAPRqx2VxVEsBWZrU4gx/bnInT7wr9wht5GxLv7CE4U4WX/r9k+RJ7FW75ZBNSqv
Lie62L9TgOHykU0ySHsvgUYYEbpUcfr80rZDV0e86WnCRS5avvTtbenKRC7e3gbbPV5nffx7HG0f
N7j2lki7yLjRi/HSID4rcpMPRocbwukLctRcvKnvKy/z79Fp1NHFUu6J9Wf/f+qZ+2Jz52BamEaX
8+ERXGBlYpUCnnr/yIgMp76l2jgkmF/nCNZuWRhe6gvphkYLdEH8Fer0TQUrmIEdarFIdveDte2S
G5qnALyNKx9Rmc5S/XED2g+jYUZAoHpIf0ciR/rHLdEg0kyK2wXExP0QDyTAdugX76U3Bbplr3Do
JvZCh+Ebhp/arhfOnwF5efNYG2FNR3ELZgE4fp6wRQ8jBalvQuBvlnpIUNDp6Lb9C5UQ8QhKZX/b
c5VKEmje3M2Scah6PrEVjbkFy+XdigM3trcQTA/nlWP3326JmNiAOvnYd5DOgHfRc5CD9uQzIqzT
LG4ssIUmc/9b2l0myBxGWGCvEuZ+/vmapglZbFtQRkPIggJv3UQMXFKfErdAFniuP64/vsoC3HiC
FGU4rzPtpK6ylxH0UpnhbydSaAkxFDSoviDActMmGr+KFk8yynenXH1h9OrJ/V7YWULLEruZ27lB
OHx78KEDlZsctwbfcq422KpbDbbKGZ9e+1BfGYDj3VUdvdFlfg/cae+T8tJusNsS6W2L6QI0dKrM
+nXNT5SURwYb+2J+RbGVOaOpDJ0AkmUpVMRjy8/lJlmwO3WB7BUEqQP36283fSgS2LK3xPg9Gyl2
O32ECtT/Z0m35FRXQ2KigNHQWBZfhOrkljmHFBQuHR0bEZTpJPvD23Xiu9jl1z/GBsVwW2cwxPWB
sfnEqV7lKmMx92X0eavicQgJdOnKxp2LjgLdlPfMRqNZFTiqHCssWYlCTbLEWLq6cM7YtydmuxrS
cabBEjQdgHgK+aOhcted0Q94mduZzn1wPmhfLuUwUucdO78vgC6Z2a0Ha7KNhNIc4EALz2mE4191
JdYFcuwo3xRh86aJ7LU+EKiHWsaU0WPP/hHMTY5sQO6sbVT7pvM7aOTmIo/IOXW1nGoUG22LPBRB
iSyMk6L2ByW6U9JvHMjI1ZvLFIhM0lXNbjZRxGQC3zvtHwbZlKZxz6DKOcscKUCydC4UQNaDiLjq
1/A9ylfGXwnzgItiz29YTBuQUUktROa7FWVHZrOgyvOZ9ebw4loZirSYKSVWtEM1D+rk9pq/WORx
HCiAfDG/pA2Ze4M+m4PO8C1oDQBVxBxc6kuL+Z0Fx01/IZ/mKv8F3AeLjQu0ruJAw4sP7+O3yXG1
b3BOKyNnx0zcq7h7dCH9RQ8sDFHmElp1UeVGQIC+Sy67p2zPq3hvPT3B+wtNGc73ewUWAUNwstf1
acMH9b4sDI5HdDn0FZpo2pvpDz5J+I1gfzwTZi4GU9X9qjieofqNhX3k0I5T+3IRc90A19X1Cw3c
4mgMWOV96Ojxff9oKwb5smxgRlSjfJp9I95u2m4zkRwgERy9vU3kRT0ZhhGNbULuH2P0dSoKKlXZ
lRer5VkF9L1LahGRNkyS/uqJAIt0RcEk/fXHXqlI5IPSb013dULUzhp+ESIBgjFMUE2NoOuJ2Bqo
5ubD8pPnFra8tj2ytC2ZpcPQaZYq1opNfFOJCkyfCcoxHD8B+3pSPJzOZ/WG7pvQG3dor4Iar3cN
8+qtjaGZWRcwW0y3Y+/LdbBSjtCzsHS2oAhE1iS15b/5MZxHrlj4FEZWC0Bb5D3gYLdJQ69esup5
d9y35KIHUcIyTFg518x1iHZgp/NDdQWsR6wPNfXZKllvf7VHWtwWRGxYM/sOko6B/bkB5DgvFlcO
vtboSDoHeTvZg5tbcMns+Ei81h1qFT+MqoPybw90bHUtmpaj/O9JAXikv2FC+Jhuj+EkvCD3rA6k
MWHGGBPHp1jaHbFZ8NYz+eophvnuHC+nSaLafHB4atYziy0HXmSvaGitadLprcfV+7RC4RWSNDuw
NPoX5Dne6Md0eFWUEDIktTDx3B0tywTj2BTv7h89mqeygAxLuol8pAj7HxuS8AP2s64O7US7gtxN
Ry9W8lAmeu7y26DpE32FErIdfNxqr2GuXbU8PB1M5/h0d5hyqlIj/iE6lc5U6QWTUEjj7+U+Op32
s+bP1HorNuAoYe20iae4khg5VEBKPeLuadKO2xfq3cFU6BjpbdOUvD3c+a0PufbqvSrnZnyHEeqv
9Zv6d9/75kgKLHM0aS9ssum9IJsDeMBefo06RU/XFvigojYZfb8iLF7TDeLymLqugYma11k5gGT8
Hp9dvnrWyD4GoIrkYggR3lckRrzexddlp4pT8fKEhMSJ89V9YzOkY25l+PZZMs0qt/8yXabqn8iI
oojSGYCMcRb3aoM7fU3Gl27loxFUAbUFOD6F9jLNpz9lE+iXO2Vx8jG1ZE8xyVWOwTMdOAoINj73
q8/TPLTDiEvAO4at54roc1xLyVHaN1qQd5MHIpp4DDB2JP+cFqzqmKMouSGq4sKD2MXjBRqgsV5Q
dt4/39boQaB8lcPuvKEziHOFAMvR+I8wZIcFq6ZeWBB2R9ASV0ltCW3UpqNKma2zCMkrEVhgFBdQ
a6OnTcCUjfymfe+vC+CjFexJVLueplIrOItxV/mnv8Y02H89kenLut4c0PHIH0S4pSX2daL3UmmA
KwVZLLKl2hmBTC49yaKy1hw1khhs8fjIWWJ0O/00va1ZjhfVkylmoA6V/MefxElOlmPFmYQCxHfV
zYr3SgltLh4TS8c+eARzrr1D2n+I/BRecZn2O3suGxlxioC0PkFnxUKfvtHxYeTi1TWJ26IOruFR
8OLnmH0lLxY+EIyYXP0VpRm9ePNmXWukMRYDbit2B0Td0foysmmwtMwkTYkO0fU04Sw29QhQwWD2
lsID2W79ofOhEMPl+Au+4pf0YDqgYZ7W2jjNfWbD8lbPkGNTkW0Vy49Hlsl+buab+ADNjsNw9iUg
wl71hRvFFbPSEMzxNIM4RgFQ7fKHWZDcjZZ+Wh6c2vrSxQXhzIZ+fXMZpxZ/7eqF6eY1d1knKSFQ
Nup0ZucdT9uxKNP6xgmY2HcG/1sgcR/d8bF7PMyR1YRohRRD5l1uElmHpK4sghO4j7JOAOn2RNrK
7DLwcBGoJyKzT3eMIpRfBedRk+3oQTaGjbz7/LvKwGrq1Kp87WXH1Hq3aRwKg1R0AFAP8eonFIky
nfG+8dAYBMQfQVSywYlEQB7ygHpE//26Vj54H9pu+ToednfDztitl4Nbem6ODy5VH7cGJMJZeRQ2
p2lLFoHRy1cSqVJEzijVFdu6TTDHg04xX8cyxG8RO4aQ4w5YQ7WkaKK32aBi2I8+5+OdBDvehHxM
bMW/PUiCuhGohysyHc9/ubJu7fixVeKvSM9V5sK/+/8vDqXlfuvsWqush+esDS5F+znBHrkey43B
tcQguw72F/0+xbzTh2hAHmTORF0Bm0/M0ZqkRDgSoA7uFpp3ya6JL21VCoBBaGu+Ep22+sYhZFSD
gNWDeXrWu9necFv1GW+T9wu1Lx+7Eoq4BNvDaEbss04FRTS5bfFli3l4lmOYdGKNFZuyWCCAGt0S
uRqXc4sEX6vc5EKq3bY8YvNGcSu5Y2nq+KeQQUnwb3qsgt3hFR7B6K7o2DEDTwI5IrdUDZW/VRXe
wYK8tVWbVXBFWfkKjpIVZLHnHveOTeX78ephuvKJN3fO5l1Pndg2N7Rpl9K7TuQdH9vW+S3fY6yo
EUhqAGMP6Db3rR6oOlk5UP+aDl9g8R/U1f/2WxiWSDhRMWmLLlNh6MRV/lgyreDmDJvg7QI2Za4s
xZyzhGCojSsiLovnV78p5RHNHQD2Y/FnI1nSxB5UJ4yje/8tFtMhaYGDyMEsFHevT2NTOFUaWU35
+mHqddeRqsOgfWYekORhSjJwfup3BVzRyNHsrtCLiEm9V3C/TpJAnRB3/MPHpuY/hhwBUDxQV+6P
SPIpjODrQkLdwcwtyTe8W7S8Fchx5zn6RyCfLWzkSZ+QRsSNCzJzzJ1/fWiqh3wP18Mnj2rL9Vkk
aHCDrKMfv+rvQOLozGH8ziZXmLuMtgEuBLD4dmlWY9Mn+NGuowsQ1x0SJGBjEJYaDaUJAsoLEDaJ
6pLKaciLEKbkP1OuxUns+d8biY9/4bEYuu+ZCYOOT8YmEtMKi4OLJH6vT+RPx/upoJyY/w36l62N
qHBB9wu5fEvW/GnaIJj7e+CESKvDaxOjlOtlBP1lyOcKr4Nj2N/AS9DdNXfzkXgNaSSWVQRZb/gV
WyGEBEfyVC9ZDGEyxRgv+F2lVgzqoMx2kztRsBhvBrqC8heyYEqjvywkIHSzGhw5a+ZwJYkBkdpj
V8lupUO5PkJNLDITbLvXurwxFoo6OdlpTwefUNezoFxj/KCXEg1eLdloXnvZ7ycUzAJTXE1ycc48
w+08e1lpNxAh8Evkm4Z5yxU5GeT3Y5ijvgTkwYIvhJzvopZ5JaK3BHjfpyolROQbx+eGjsP4g8yE
xHQ8beCiq8o03v1GZVDTw9NxrzBmiad9jDInd+VyIx8SMF2Cj6PkoG9/KnxUZpzWYZG+L9/I9qZc
jrctPYcXMam4yvaj547m3b5QnSLGelNOXLqBd3eAYcohFNwepWmyPpyILqC/uhbsAG05AZKU1DkJ
9QcQwwgM/EqyeUUsq59fVDDVmSw4SZP+odOn5L23lYF96TetglbqbMb+GJtu2BZn/En6hoUiolZI
4ruwkRjmkCrsZJAKJPbMbSeRJSr18waZbc6DCjm+NbtUL3PFHlJb8I6R6zPs02Q+9WPy8ESUMFTV
+8r4htjCWS/TqdwYWYKqdLRdHByKfKuNgN4db57syC5FHV7lWHeC8+ipvobQE8GYsyw+4XUIYZrZ
eKENqTbMAuvECGY4RnXCJOX68GwhOSkpvUMOstxyCNvtIwWYxbpOXObN3noRVbthwrX1qvbfpLib
BbWnYLZ3rpijz30YHN6vm4OlOZzfZtE2ixdBgp+VsFaAMiueG2Pa8vqvy0NRHPeOtEuOn9Gbx2F/
33jnwNSkM2p1sZSjuJw1M8swnr094gEyC+gHf2yO3ENxKZ7SB+mn65jPFL3XrC0u8lHRsyC2Ekw8
v2CSXxZXMNaEWoAkHhA7Ws+v+AkRTJ43DebB9y/X1zIpi1blpQfsI0WQsIwMc7cjHF0JHaN21hQS
t5ouVNhVDY97c5BbplT7M2Ne1zAetniSb6VHS38sCPr/GvV4xcesQ1E8A3ztrY1OmFWAGZqK3uef
t954YmggwZ4VqHwN3VRQUuk1RoEqVqNGvJdnuyfq80a3CFmL+Mjg2Ivb5/SXADU8mTFNtez8/u2U
41otcP+RLFoWYIn1SSJTsrEqloGqdHdYULQWKq3ODxn5Qau9nUHJ9h5OMRtE4mE1hRxo7lNLxo+Q
gUlt97j5tRhZT4exhuTKV1QM9gYSAGXqBLPgBWBhGLXVFXLgUlwdDMpcrmyi80FIvK8jDo/YmQ3P
6uHPvszHHHMCQEjTZyx2B7D8d4O1jsAcvYUyp12eIWLiHBw4KRRLdCkbW6a+zdweSGq3De6/qTNM
XWpiX0pTmDlsMWvH5T4cdLVwcmp+dsvzaGq1yXaCPwTnQZChUo+M7M2bRI+KNMC7MLMmMIv6zmhQ
abzB79ZGmARJOtR0KmiMZC+RezB1mLgVEAzrXjpjf5uzdTiYzcBX0q5e3cl103/o8VDyGSpnW1qw
5b3JoedymvYcgRvSz2dWanx2zwTGm7KXij0UPp2SsxNdkNJJRf8UD9rR1z5CxYzhcj/TmgLlzpjn
inRROiKIDjk5kabK+ny8QIv12jMl6VT8ouXQLQC9UVQB6sLP7BebrCPpfJsTRs3mzPVHfgzRtUEo
llOSEr8RKYSSFpAkuvKw80bYhwRoIXZqbY3e3DtBYut+JnZ9hNJta+1S7h7Thdj3zHVDn1XCUfVJ
WsXc0y22tvKXBFIhDKpgf3hlCoguW6ZUdS/Wi6wEThA+dYe0RvepHjOOB5e4jHGb1DH+GtTWQdUh
nkRmXmZhN6kMFlHSxGrBsSFrHhXORE5yMKix+2v3yC8dmXh9g53GGlduo08Y3UaQmOnR5AjNEGKd
oJi7WRLreoHvU+IUFw9GzLxwTVjVesj13nHhC4lzdg7zvZQcAgXvckD/GfKVgn9D9srkIaaipRtp
QMFLu3slcbpb4OBJvSlmaeMbNJOOwZN75iOAQONcOtI5H+RCBS4jP0b7G5AxvfeqG/XxzJldGGdJ
erx53gioEtxjgfkE4zEvdVrWTtx04aLEJjab/itrQ3/03/w4SFuUkzwJTkeg1pe9lXac09JLSfR5
MSze5nY5TuQ8X9eVJG4ysX5NeO7+/qrnteesUDzs4sbR/kxRHqX7lypngzA82NdH6nTJzqkKeQQr
SU6CxHT+OpN3+hMdUVhYBpeNTflOd70qHRQhxpkV1DSicBUjOcy69tegO/CePPQO5Q5ptOUbk3YU
fo/yE054Sj7bnKRh2XzWksIQUMW/dtPphUYW7VujSddfJZQbrXxT5KfaPuLukFovA4KETOOebeqP
wwNQ+xFdWvIXWhTMLxDiJuCKwPuLawL2D1OTgaXSIS13rS3KreRovfV1HH6C2jdQmdv0cyM+l4bV
rxQ2kxh9EYxoWdVqLjThWkrYGs9ECqmoDwj1tPtJQscuxuM71Pz1HLd1D20YOdfqA+p4+WKTEwZK
yXDQ8v3JNLAm0ag6/pQNRpg0iy8DlcQDN5gqM4Fj9PEY4HbmSOHYzF1Agl8YWAgi695bSBItqV2V
roT1n5T9eZdXfusVZ3+eJcJcDPLODnU60PRyPs97YyfEBxdfDQEAh/qVaOUX6bE1MVDdMIhVGm+G
lyXhvc5HBqIYhGCgeOwXRai1cIX+rb0pD5Lmmd/IB7hwkKq1kFhIjYntQBnUG6IMBPv+7FU3L0iV
b3rKfRZ0GqmO3p47D6nwcSB3fm/NdRrsKs+tnLs84M35upbp8r6cKmmPYqa3yR5te4uhWUS5yrfn
qKfmu2kWYi90z+Ag6gZQMp3oWQBcGhYFyjSnG5qUOTV0LE1Rsk3n1K5sr7gdzRrYRTY6XHBpSDhj
N8uD+b3/frp1Fkv+a+mmItCJ3lYfiH1CBuwMy0Na1iHwWJVeY59bPen29mvPUpCtruBJJmr+CH2h
tx1vzYi1pBmKnxd3rCZ6iQooBvhnIFbhS9s7UWJxgwHk/rdOAjQq73+TwTMtUv3LSIMgQwJBL4c+
iiSHMrvdyB/XpT5EDTE3y04VtiP7f2bhBt0A+3Ol12lAvxc17LcbEbOXFQRP2kS4igC0v8PCpr2E
V+gmNIyunO7v9CFMcpuU+vVO0wtEvL1uRIcdnF2FdhTnZz0KHzdnFUzVEi929pHIbF+0gr2v2nBF
046YMaiTn4B14nZ4Cnz0B9En6oPBe+uISf9dNmoTXr4uE9ga6o0gH0aVGCZRtvIcuoUI7KDh4BHW
RWYOmy7TWi4qWZWlROh8gMAt35WuJ8hdYcZAiw0IYseHoC2KFBqSfMbjoElXT0p5UZS63/Hjpdt8
zf3Aq1YB8cMkfUXJeGsuLroJmrJAJtReiEOTAwgiPTr8Lu9Ir34BQGBwxNI8ZL+R67R/b7F8kG+f
OebNlvmDrx1TsCBKeVjkbYQexJ3QkuD9r6W9fcZS4k1TweK8egYoq5fkPEx66qULuCKJcf5Kk6Uj
2yuEZxqMVoEJM8MSBtyekB+qu7wJ4mmUy4XN4BQbNFN2kfwgHdsR87d90G5+sDecMT63hTflPppp
Zig4EEvtFj1+fo6zFebDr1Wy5bSlGT58l6DpAUd4rlOQzytCS3TQNmMuZu3dM95cwNWicIHw/OBA
qvd5c7s799Pq/+SiLXKKa5H0yh8FyEDcTWie6ZCMr8qlU/KDj5DHdwfGciQpItqa6mjobcyBWyHR
2IoNVGOKnIuNDZPDX5b1pYXogy7cInFC0oCGws+vBKKeboPQjtTruGZOOaolXNXGl594vBvfLJnI
A4R0ezUH1XWVwFPh0BglmXDHlKIU9yAJLbmI5xsHscOA/1PS0p2ddXer6comRmvTDDa04830WudJ
FwR3uvcO0jD5SlwOqv8oYVkBxOKvjxs2DIV0Wo8IGM6rjfIznPJHh7mVljaxz0Svml9lCTroDVA+
s1x7gL4hKZN93KQSwC/ou97GVdLjHKDknvtZyT2Gn17yjr7sDZKZr+JvLiOqfnT9cVnbDTLUvODu
VNDGo8ImJ2ubLjTK+/bVz6iP4WFk3dgLU12rG7TbYEAmLV9ShOMZiMDASsqO8tnoq/Lkvleo7tdC
PPe7CDlvbW9lHyM3zf0TW0YEcqkWZimznQqd09hdUK27S3qFUA/jKwcBrcLcsr57no3EvIol0O8b
TbxQXVLz6+gJZxMXYy6fAaN8IepuxFl3qnux7dLkmI7GJWvb7iy5qNDqonP+qu/mDtvFDxECaY/I
/6Q8/EPXGs5+RAeigFilptXzjHJ3j7lYsc6qoZ+BjQkDhj4+sxSY31YiIV0UPD/m+6yQGMv4Ar/7
DkEMaiNE03c+i2zLLJKzC46xaPAVgzq9NO1vB9KsRQhHedun2Aqc9RW9eFfuu/XmMMe0MVCB1sVp
HLcNbgGVJN4jcdBtqzUJJWQqBqMcwqodVvrU6jlLS+XtWZgAS3mlTcHiZZTn4B07WjtwR0XqHHI4
Tv/QNnBPZzUQ0cO6ZfFNRyi4T8rHcJgUAtrq6/A4/JgPM/wB1tIY9OSaxNfcz59zeuAHUbounNKR
k47XSKTNCHHWs3mNhtQGed+g01eGndOlT2jUhocGL5R7lu9zJCatFK5YttkK4xRrk90FAjCHia8V
BDRHYeGpl+sLEmz3gN5/fCd1r8FhKWnxlC9fbsMWPgfJs9lOSK1KoXL5HvLFEEt8hYHW7HomveAT
x7fYfBeQ126buQQADteL02s3VoiYMC3/WlfOw0h/Yf7u0EjfuDSbNBdEdwC+HvCa038ccC5LszlH
4qJwxLQ4zcXfxFph3+dLbbtIsXikLml9vDL7WyFFYyBq1p0fPZRL0ug5U0ZIjKbZuHtMlJ7eB/La
6/hBmCoJrrJP4iYF0DOYjtJeEQBy0tbF6D3MnVdv2VPtN72XDOzbO0d/VFtJ1QcSrga492mO/sSS
zkkncv7SSW1YtH77sSMYyrIlerCqgF+zm2JzXncl8xdCe5jhRKa4LZXRwUTFSoxkZiC5QncY5yfc
5+3d7qMw+te+bNQmKrSsW6pG07c706CuNwyFsjs9nL+ws3rprChHfVw7oui0wDenr3ukaxmaS2uV
eLtXvEgiuEjda1eEtqbfQapnayofmYtG30LmhVMYjgOeAxY2gvS8b2Y+5rPQiLsVt3z9Xn7SF8S4
0qqblCv089jEQ/FIbcpWkiHnf3Hcvdt+82jD4YvjmiGmYD/FsvqCZz5kjrGU4HmLL6eYRmaXo0wF
I3qxsNfm+wWnNgy5ghweKkhUZ5QmSCcAsYsraB7ttojE3do5pBbxmJNCDSSLhXZU98aw+/Oc8GCk
jWmBDXOdZuR6PKg2qwW7RCr808/ePWudtvEd3nT1SBiDxSBaQLZXEqPN07R7yABsviodq2crXkWO
vlkuCkZaRgUxR790TOaR/TSiUazn/3DE/39Pzw/1uKLdXGWHq7r99FeZLH2v6tl90ImEu4KyPbCY
kxvcf8g6kUIiBli4PDycqeOPxT+eL6M1c1/YCtnrOi9lBg9GjFsDesszTL3NM6KypCdKmRXgE6Gp
2Rrc9HdL4aVypsubPYrMhA8rCZYS60m5k26DGK5WRogA/He9wC9w6BGq3MatylmIxoFMKFclFSu0
+qamoyPjWMR5XbGetUxyFTykqzKS1JAik5p+3kQuZt+dpig6u8A/Gm8iX4zJdZIMGXXnkce/4MQI
mAT31IfmvwwyC1HiIzKFRJQCBp4OPqaL+qXgQipn5Y9LnM4lXg4bgdioQ0iuWi727IF3OZIGUvAP
kJcL78RmiEwnDiwOupRGLIBsDygGoyI89Jdb8bf53dMTebuSBztHNjowhJeYoH6ouHvW7R67u/qV
pOJUIt/hKI6fM8VLfdLAMHdcHy4po2PVqMACl6xPeuQ+RfTMo+C33nLrv+vHCVRdJiEKwd6Et4Ro
EDgYdMc+HBJm9qpxCsFfeinyKS8R7RgRVmcPbes7C23IDdbDkh36rZXLBZ9Xn7Ow7z9BV2/NMWjy
SCzOqMGzPROX7h8rCisHjcbqm9fzX2QzsBx3w7RmPI2adcPRz3R1FwlkvJEHCU76NNDtr1htoloK
5+IZFnYxN719L0qRYcoSt70ew9VVzPFiKb7tQY2ayTCnnUbwxEzNWe2LqYo8TfPRvaxAd5JdgaGO
g+M0o6HUYBs92iplz+iPcuNHd5+vnDLSejw6OWV4nBLXrxAs0Hnz32QU9wS56xnlRyHgeVQPM9Gz
i8P1G/05WQbYlHxUeQ3+GcE14dswNIal7yOwV/qfb6LdduRLdFqBJy45FPlecVN17Y/yrmp+bo38
gGRX5JWXVORIOouwEnWJ0YYrR7b2IAwhlNZvoSCGZg7BUMIXIktTyKWQhDzoTuvjIC5li0pPVJ+Z
EpEsbIyMuUsAFqeAjhagm7aRj1zYXyb+etP8Fen/WeJCovOdK8ZsxNqsZDpJXBRJ5lFQMyfM4VFV
kYuAmqkaFPm/7zUsN6N/KY8cpQA8O8hFfd1f6xrqr3iMaq/TFJuS0yX4B6a56droC4IfS4Al4L0K
WgqudsUfF3kdUX+Q7hJZs4wSu01nAtio2T2OjqzhCY15Aw2HwsBYUnssS4eVBjv+TXlHeqD8y5iX
/a+lV9sxMJF5tDFIufJJReTa2MT7C+VJyFLT+L8qWAwgRczNm12fcaW5RIpUNdzYuUYbeqdIdd3O
78H+Yeiw0gUCrqsAREOtw507oaZ1muylVNPxTuKhCorMJUVXQkVF1Eji2vXEe7mBQsYPZnLg9LfL
D3UwtPcL3rRD8u3pr53wLVmcJfnTNBaWirsJ+Iwgiw/QHojbAo2ZzrSZDJFogsGNJ809i0XYJJ2k
zzjBzCL+MTOjRlvURIB/TMI6AGvEh5JB0sU6
`pragma protect end_protected
