`define getname(oriName,tmodule_name) \~oriName.tmodule_name  
