`define APB_BUS
`define ADDR_WIDTH 16
`define DATA_WIDTH 32
`define TIMEOUT 16
`define BPS 87
`define IF0
`define IF1
`define IF2
`define IF0_ADDR_START 16'h0000
`define IF0_ADDR_END 16'h00FF
`define IF1_ADDR_START 16'h0100
`define IF1_ADDR_END 16'h01FF
`define IF2_ADDR_START 16'h0200
`define IF2_ADDR_END 16'h02FF
`define IF3_ADDR_START 16'h0300
`define IF3_ADDR_END 16'h03FF
`define IF4_ADDR_START 16'h0400
`define IF4_ADDR_END 16'h04FF
`define IF5_ADDR_START 16'h0500
`define IF5_ADDR_END 16'h05FF
`define IF6_ADDR_START 16'h0600
`define IF6_ADDR_END 16'h06FF
`define IF7_ADDR_START 16'h0700
`define IF7_ADDR_END 16'h07FF
`define IF8_ADDR_START 16'h0800
`define IF8_ADDR_END 16'h08FF
`define IF9_ADDR_START 16'h0900
`define IF9_ADDR_END 16'h09FF
`define IF10_ADDR_START 16'h0A00
`define IF10_ADDR_END 16'h0AFF
`define IF11_ADDR_START 16'h0B00
`define IF11_ADDR_END 16'h0BFF
`define IF12_ADDR_START 16'h0C00
`define IF12_ADDR_END 16'h0CFF
`define IF13_ADDR_START 16'h0D00
`define IF13_ADDR_END 16'h0DFF
`define IF14_ADDR_START 16'h0E00
`define IF14_ADDR_END 16'h0EFF
`define IF15_ADDR_START 16'h0F00
`define IF15_ADDR_END 16'h0FFF
