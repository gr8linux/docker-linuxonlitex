`ifndef DEFINE_VH
`define DEFINE_VH
`define module_name can_top
`define REG
`endif
