`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
rODoOdoVwcZ9YEaNHkTpBu9/eCvGEoHnz7UkhWktIIQCNti0dSD91Rl3kLPdL6bSdvejXB8aPuUz
67UflIy3W9m+OfMIMTAd62+bQskPrUSRQugufBmEzb/TeBL3FcphooDx/sflJfJeTvXjRF8IaONX
QakUoEzsMZI74FO26vkgzkXD3JTsJ2u5xGK7huowxWQzowde11qZGRhwqIR3Az0jV+3QLxF/Es3F
RBp4Dk5KfpmiceJr/jzBC3ufzkjBTyPICY7UrD8eXyx3DRJmyHU9hMmuJj2FJIIlZ7Qq6vx3sGMy
yytNlAQbJ7McAkU0HqusvEffjBr9qnbwCSrkaw==

`protect encoding=(enctype="base64", line_length=76, bytes=110752)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
UVwUn0eG0z/fBvABIiNmNIfpBHbzDdiHaRbfvLyupJJKNa+bbWrjV54teZ8cSgj++IRoHb71LPcW
ovwG9Ec/g7dgfijUQLAGYJEP6apmQoomCHJgBv2L0vwbm+lk9sav56kiCbNDY7o1DA8cA3uxFT/r
xF8awwkr8cG66xb4j7tPsuDRsb5P7aoAwTPOLaL0MEIkQwOqrJwFTzqbQ8lfDSX4Nho+Og5P37/n
WDbp04LRYe9CljuRfbWH29QfdqsQl7HEzBdqzrWyDuZHTbV7tXlZ+YbCGS5r1JVud60hgllbLYI5
PTulbD/bHe9GpKDM/1H1pKwUGYJ4tQIB3bthICPzqWsQpeRpuwjB6RENaFL58I0Jr8/JRmdKFKM/
hWx0e6v7ixbyjk4Dp0VmqsEu8sRCSJBn552zf9KUeTW59Xb3QMGz+iYbn9YZ9K22vGbsQ025JV33
20vnko/3IEjL3GEEVNAeWZERRHJLArP6TNgY+y2Ygwvr1YI7vK9kis+PgCRN2xqDlBrpX0c+Uuf5
BgyohWIDl8TOG5t9Tb3OZBLrx1PeS0EVsCUge2+PW/ZZH9Hynzhsl7EayNCrpjL1hXBjBx2I8Ql3
FwA813t1vvw1Z0zJIsSoPn5gxEcPEkNrzYNkB/8XQI50eQWg2s7o0wO2iM5nvzMexoEx44HzvTfi
Jm/FQuop9oT5Wse0fQb2Eopu7fclcI7DSjuZaXNOYSPH8KVTvDCkpl3vLHWEA2LyblNoSoaxGedy
NcK5VH5bi8B69TO+OUzY+5d7oq81TaDBy3rE113rgbNAp8NulzGe+XdiHGc87C+ZgsQlgsI9aoJ6
nBRrAfQHQ3nDABNce0H2byJv1e2gERs+0mu/CUN1HcWI5Nyzs9zHU7irZRNYmgTOQqg58aQ0lmdP
WkOOb/pDvs4mq2TwQGanLwcwKBpsbC+/1Hwv6vr89tbNFFHlL8fFaHNXBUM7M8ahLDjJ7I5QP6YG
XOeobh+H9X7I0VorQkRZPKm3jJhG5xai0lcuh/Lj5EeRTJKnQUwmN0DWYSYbM4QPbe9Qt10kJdE5
qHKr8KN4DMJHqhavNP7L1EQ4sIw/xDTwNDh8Mb+czTyG+Np7VF+1U1jSLmhZ0uC3Bh+Dlm6IW5ao
pTxAGFVmTuqgTYBI4zcScucxtW00AkR3aAd5r/1gp11wGiXIjUcgs1G3uTfmtzSMFBMr+2liAFIh
MwNmI3Vqsos5ecEc8KZyQKeYNjNz36TFN3aQjF2rw735DxfJvXjtbIEgHeWdQcsb2Sv/tTy2qJ85
6UUWCINMwq8CvatQMoRFpwdl99QRQpAPXv7mvSBn0/8+PD+eVwA/6bGH5SDjJ78IJv0qPqRQwZAL
BgEcHQ0iju6vZxru4kr/4LxU74CXnxfs7OMOAGYRwRKk5lgkLEw5vildzVBmLciP3mm8993K2ToD
fdteP3UPNLW3WC9Q1nxADhNOHdzlfDrZQT+/6N4vRxUWEJy47sO4jWnDIIuJHzNNjKZTU1HUuvcr
TIxurWggvECCdcm2qYclTeU2yyho/5lSznpPR8o3KL0jMM5HKS+iZEl+ygrnXl0UTvkAmWp5iepp
cKSI4qhTaQEVz7VYfGE4oyWE1ueAy0m954/1ceAqOVkxtuuXbIhw6GT2Nxr35H+iu/Glm8t03pGG
z7a1bpfh56Sml0fb1rsjG6SsKnMAkL0YBuvCecNyHw6F4CUDXHmsvMbbzkzVmOXApNl1fVclGepK
+H1C4M9OgxliwtATdvaovDTrxTR1tjdJeigE0z8Oni3nTzs7OdhyZPCK6uCwbJZ/CowndofXPoWo
nYwVpirkZs1nh8OxMRcSUgDdxKB+vq8jPWGZNz9YW78wrOpQIaSinBsKb4jVTBi0MAnmWvEQE6VQ
Xv0pXZ67WZvfm13/+Vgi82hWPBi5CyB3kB63Gn6gl3HHM+yqvQRgQTPMlUtpJ9wPd3b8hPzEmFTI
OsYnAwlQjdBz78pETJHznMUZY9jFDC1OUkvTfJj+IwJlKmhq+OUrf50gxQiX27YWTIUme5Gd6Eex
ujCRe4cQxTZ37m9ezV+UKEv2l6sjqH/iC0DnoookQ/nzSbhuby13GOH5H32W9jT/ajIOIZuT3HUO
/DlpWLYo8iT6aXaqv0eh2motzEyx2lsS9NPeyJKi8YktmUUtWyRTUdjFqEhyZzgpBlP7iAjCMd9F
W72xmvpgN2tmxLqtc5fPD2ONgfzg8At+wpvR7iSIA8l7Tl+w/sU0dcxiCeLlNI8Fc+jjuSRFQitA
gNQCp0897WBldSEXrf8IZ/na+qyPnSTxZ7CTfxSOanpOsmJdRjgp7/1zCUPA6FEnvCZg2euIk9r/
bOKk/oKzM9i+OR2iS3GI4Gkn0VL9+Sh789AhA54QslOQOMkoAjPAzeKxyJeotNUTNBVDl3wlgyRI
At1VXrXtzG/J8Q8jpBtVHP6zPd+lAqRNUFH8H+IbaUSB8tMRqrXmeumlNSLZMcbSSmFhjs5N5+bL
JPo+Gpuv3oWUexfh68h4Glti0BLZDc/aCSOYBgJx4cedauIloJ0CtZFin/+PGG5EAM7W/Hr30NOh
dSoXjX8euEsWQOvkNkbHGREvWx5tyVTvwbr1B8qeSO4cvYK/1RL7i6T7Lu2330vwSJcNtE1ws6df
mWjI4EWDSpX0xq+bTpNOJVUHTdR2jfrG2lte9n8qHZim6enJSKGDXj8SsUahhv5l9a9O1Erp1F2X
otTXQJqWGc3wDkfka/Y5S0IhcO5YFXUrkfRnSod4eApye1SPFZFkRwbfncEaUPMMel+iw+7mBGI7
9Ag7q+EjM5NrPrmD3bewShY2urdIqWkxzdZzI+OE1V8HKKZs1RnMZRTpZmHbToLUFSAJljwNJTXX
UPhmxvqcsgiwu2q6LgH6LKG4fp/0LYk0AcuYIfLIPnQXocv9iFrIwmE/7LpzjbCv9tLoiU/qX6QK
P5px9MltlAnAX/Z68kaIvw/NH3AT6K6VV/iljGBg3+f0nOdwkPi9RLjzbYqcMxt5visPosn05s8R
BizECearK1MbTigFQ457iqTYrjaOBnKnG78t3Mk+kt94sM5/LLfCsSwvN/rPbjLVlcaNizHmqO6y
dMQjlYW79aX2GII6jz1Y46DIjoFOlufQVHVKOpkAv4/INXLTen4+t2r1MSRoU0sPrF6AM5miJ5KU
75ekLow53haxRaGU50ozWC8Yapw4AJegMgt93hn4/JFkKGq9Vm8dURW+ASFNaoRgdW2H281DNQ/A
wdt3kFlsDe0gJi17F9QMENJIgdZlpq5S80/qa8wquKkQh5QeMUdPIdyr7R2Ofa3qD8t1J9AniL/Y
tmHOSD6fPgyYOhgSNUnq4Mj96jIiuBi1SwpBFdvzHV+uKzTj6VkLXjeyqZNJqOvhSK4S0HBrU5bg
Izc+nt695LUJy4u4YY8tPZIX9mta0Lgefm6WGlhrAUgk2COAo3I4ysnWOP7tY7BqL6Ib/8MDUJ4d
BgxAnCOI7ENylT2RbY72iEhECLlBjJHhqEgBXNVLzz+PrMYP7yaKvw+RlOvn8K0Nx99igVR/MEAF
R795dDNuJVF06R0SQyEPf60cXAe+HZdcQS7E6MtzqNvM6V+LgRC8I0ZX5yfnCf1DqnWHKaQ8+VqX
0+O3B/0IwNIZJNVqyDI1FTUfxn8m1yet3vHBSTw9BVOKooJLHz5TOFCBre2wAgEOoECKxsQlgzpr
UrXrv7fzVdx4turKyAQ4VyF2XFxfY0RzE9ssayKerbrDrhl8Bx7BINNbNkbEVNSu1s1cQa074sFX
8gI9al99pFaV2FNwqHxtQ9C8iH72DIuzbjzSuquj9QizQ3M3XcrDdQhLpWl/bIZ0v0C6EZiN0Vxp
UdIxs+Xpravn/yavqKAQSZT20BeCGcViIaBDOVQqsxa/4TeF+okKY0RFMzO2M0UgXK3/EwxoiggR
M8guA/L4OWdWWcgkNiszoWzdnhiFmEG7UXqv/FtX/Buc+JgtyJYnb5y3Lb73eA+YAROonTFUe6MR
Z3b4JAf3eLE6KHHmol1rU3XyYZbleLw4WifaE8ek3lF7QikKCfg1yAgAylb7725lzoUkMFXmDzdS
juy5bp4G3h1/AIy265KTF3ZcY5l5gQ6p4AhXV/5fWSI5Q+cgTb9CVFg0T56icSGCISsOMdrvr3Nn
Xinaw8xhb52ZyQ12se+Odaih91+1AY40Cq18w3r9u6RNEPSq+uElA01vI9HK+KPSvBdgnpguc+/7
TpDxgOh83xhnf6OMRFRpy7BdGTK6/jr6YWg89nBTTBBRijEQCfi8z3+DUPG964zi0/zI7F3+5NeA
lKACsLwmWqdwxM0uYCsocNAzSrIxzYxNRs0NRsTf807EWfPIWkXMFV87PCKbFflluhSB5dKNNCGp
HFoYUMZqRxzxLfZ2bRp2OA3oa+MTJlQItWQZruFaJTc8bfekA76fy+BxDk9HhX8GsVo58/Y57zqr
KbA52Cxj8TgeHMXx5jQvpmNIyyxR45XnKjADz7w8ZI6GuM2mylUvCmlcMRhKLoLXk0Poy3+PkaGb
VjULCPrhpIBzXOANHUQ5Ru7HgpQ33ICVeusduvmGr7mlaIp4J1dSzwp3jQoy/ae/nefhg4fjHGH1
Ne5oqD8+6klDv0ucS5/HfRfTv4GDTvuAxCh4Mi1yYi3ZAjGkQfjiJ+jRTBuLYaL1Y5qoIeJRvTNK
wge5fJb+/JjpvJG5sFg6naS7ytDgeBL+0eLb8hXnnPSNGOhw2Kn1fU3GqOcrd6BEV4yPPxCLMfdo
tW9yGHMILBk15mcPCcFsc/UBlV/rdQDMREVRJ6V1Fqoof/sylK+66yTK5Lzpe7Z481pwiWun3xRP
FW4SZ2W2XmL4QgLTnYtbNjX5I1RNpfXjjtlN+kVaQCKl6u+n/3lMxzUPrFJMzTDuiTyczbq26KxD
6VJ2f1X549GlVsHwj68sod3zRgg7RO+6qFgpHuha0SQeqKeaO6VJCpatM0za2j1UzAxeprw4mj+8
FrMCAJVH9U4OiBZG5tLVx4qcAIPL4w/LXutcNHtf9vX7cSCQVGgk6X4UXX9L+0I6O8+YFv8/+SXv
txiCEH41U2u+lNBh49m/S80RZSolTcBAtth1SPPKUnP69VVqqT62Qhmu+0i8hBuR05GQBO+HsIxM
CPPnkc8QqUjSFcniOIHnhhneojzHM4Kowf40Kl5upT+2se36Df1VhnW+KJP9vqHzUUlCkH3I9uM7
jU0tR+UccyOnFbaQ0FDnQ4b0x9xgO/dOk+SXKjVts4HJkdHF+ewSy6ICuvdKbVRx1xCij4cMiXVH
f/Qrhu19dAjh3e2r8JTdyyGnaiK39JLjSRff8VBz6KDXZEk7/uuUoRdxmGOlRRXflX8jzvs5TDym
87Djk1QrXl1HIK2rMdHLLDohXwP1ag7xlrnJNFnI4Ma3KRgGIp3zyurX/m0YH0Uvqg40EP7r1jL8
UjmfoCU9qiCi7E/+PqyQ68gMFJPFSvVvw/KUe+9Gigno3u9/l5xjwEi7FYsKZHiL0XQfSyS+pOvl
eGo/gHa4oZGdT6v/QE5nugm4niQ8+ZSRqZVqyaaCLsclxFm+Qv2gzMAY4zBqHKgsZEVvecF2hNLz
XTPhQcD2Y0bIJmO87QHOC4SDmjhkntTvaIZ32axuZkbLo84Hj5NacabmsX+/hohRULzjyQYhrzJ4
V0Fsel/mE++np2HBh4wTX7xkrLiB71YlAICGuKzVfQQ3QXDVct/XajgcRQUtCFR1Dym/E3lrXJTG
fsirS+i1Qtsrq3xwJyn+2ZGpcQXUid/3dL1HalmWtMi8f5DtGAumKkQFhLtzLJyPvDtoX6YNHNJx
z7yzqwft0Df4az3utvpgvN6+kMFg00rZXuaAHcQmVIRGnfT7dGyY7V8wEscEOAExT5PbLluo8agi
ce7UcKgrH/PWFZWYtZXrx3T5X+s6ytv1Yf+xeC23J3pMzzmdcMUroAM4a36tHd2g00tfwxRqSaBE
C0sdRcETYX3uF8gXM+RaSAHZ3pFH/Kc+Zf46Wj1QcA+l0DDzR3QLsPYD1alAGILQ5Xpyifa9Rt+T
zMb7lTyb3LzizshzE63uEY6VImm059TLvQgCRFFTejzIbwxIwR+Q09hCpEO+t7HvrwJtYETzY8vx
J19IhK9QJaQ6w5AiW8pN0SQijTs/XKsELbqrbgGZ+wL81cDoTssuI+ZN8+/4vi+D6pyAsrr7t16B
DgCUTGWrNTuokb3uTdyhqHVc0NYHHh3holfkwRCDt2rcchpdrlrUPjc+psVGB4BfB4hHbIEiFvlD
xS+Fkj1/W+zD+WQMGKjQy/v2CnhfU2C5WKyd+0km+Rw7G7fn85cvnRUOTFCaDrCMB8BTCItb2tja
tDbApmhKB/lRhiojujqH3HcvnqV5OyrHjJ+oY9lT1f5UeMU7RLnbXTojMReYnadXJ1mm3iINiXqH
ULbsw/ouVGV7OmAb988xP4DGE6PBynkx5WS+b8WyQAZY+dRraBbhaIBVhuqcODCfEkeGw8ud15u7
x9oCwPFTY5akX8MIcTUufTg8fKFq2HXVW3wshsd6fi9R6dJnMElP7jc/M34EugexaLkkABn6ypsd
xwAdZlX9nlt5VhrUphM1HY5HQLh/235dyfKcyvXO3rhSRHNTwXJrYYtis4GOrzyVlx/hzYuaUEAZ
+ABEKmjKlWMZa+LoEhl3TENlTxk5Y6bto8r0nGYebNgLqkpNJQE18RQBdb8Eky9YT94Gqe93cJZa
71/uiJwyDo4VxEWAb7wsqMh5J6pOzo9M1YCE92tqCmhW4KXSbzCHHUwkaxLfrLX4B6HbjWRqE9Hh
RQB3+5oMm9wgiHlZF6iD1Wl4O/NKb9EGIsWFzSRWq6+WDNMRqBFaHN3euSq1rJSYlm9T8SgaiXVF
zHLUO2foNlAmBMpFDG5/ERasjyeVy5Ea5mX4MEedIchwSHraznJDeM9dsnrkk2S8TjMm7j3jq8Br
Hmm7khFEl52hrOXcJa1sruWWOJqXpfpsjM2mb3fCwND/Q1cA4gWTQaLVePNSLMThZWDRyNp4Hx3c
ntiNORv6sRGyFaAycsA61z1Cne4zjHW55cVDxsgt+nshg/QE3G0oH4HFmKzeVwk6rRtEvqrbcMiH
O5Nd4FiRxuRRFlHrKjdM94txlnTEDfSI7YBN8tyMpBlfy61hnu1RsApwjx7L7JIJfbKRYMDwvyrO
Uo1ix3muzk0WeKlrvVZojVHYgRRrK/J6M0EJ3cu+9dELQwn6rWp+1q/WMPtTVJNho31ExnG6Zby3
vB9Kxg6khMipabfIF07FpUowHNf4KTxpPLQRBa3tSFGiHsZ2S1/RMsjFaRY8bFGsfhXUf2CjF02n
7/6ifgNHyHkvHYr/uzkmrfEIt1oFCfn/g2HSOBuTOoDfX+M13quT7zSP/LqEBJznSvgAJWHbEJeF
Ll16m2ikjOw1vkntZ8rNlJUm4JotGNSM/EiW39+Thj6tR/AaLrWZ/bHO11Y4L5yF2c0T/2MrSvdx
cwJlo5dXKY6JiENEkaV14K8sjc3pduZxicqXQ2niU06u0WcPAaVU03sLWnXDpt6fLN6Xr9fA3ETR
aI8ZMdyA0EujegHe/+BWSHvj8oRw9j4CfmhLmeuNQbnOJUSpYqPHVQj4k+iLVOraQIRpIEi0bw3j
lfzQ6dIi9bNfDLhzK99JJeMXefoKo+Gkp4/RBnP3TQ2wC+qSBWyrd/DjCOCeH4xzXvt9TfWCckT5
sIxYADO0wiy1eOa71S3PXwVbcHkEGUpP3Tb6NL80SYWnmWVrRnEwFGYOcGPTWObS76+Qqfy8LXn0
7S70bnL6y+GPspPS4ZjlxpjTvdWkoD94ocwJq8ByUpHQRm4xjFeW6PNJrm0Kj2lKL8HmobaanMSy
XgRVdlLFMJnE68mcPEgAZn043IbzgkttSgj9gqDgGtbLOQ0Y2ppGoNAf9jBniJv+A/3b8HMWv3iB
olO19K8On54itd5x4VbZl9RFsGDE4GOkOMw4kQUG7BDFxYqgiV6+k8wKKK+34vTX7sFObnZ3ij3J
sYxGV0/7W1yYKxCkexo5rdpQycLIc7tDkclmIbLnQgfU0RwKUhtCTHzK82zaMZO1ur1UZaJlLzPS
xwVkgbQNUQgMOMHAWWC9qJdu0QHBdmbOFf/PWBJDXAhn2++/sUH3cgcCVJRI4LhjSZlB0rFRIw0f
p2Lrdt/tifJDssY+GCPvZa35C2j7m2xRPw7dRCb6tvCMx+dnhIKN4pAzvy+amVP9gXI1aOVoiytA
qbNWX1EhQag5fDDHzxNdEw5VSfpXwTzmldTnGg+D8l2AP2rZ/HBOlR7Dcng296W01sMAfN4S6Itg
ycwPp35jC/GlM2fuLuhDkVzKtzoTBQQwzA+LXBTCmsjSUz2z9XCF5/BkBbR4cOEAlIw0vghqPGP1
fpWKMKUX9+sSld5R4wj7TAZqNSgsimazsor7hNgdejzLpSDzuWTqHlFfta8RcAr//CfGm1NeyEcQ
IdLzKjK7zOvQUGosayySaQr8386bxtsnS+Xa8QlNF416zr1MoyCOlhsRMp457eaf8Cfg+iOm20X4
Jr6bzQk9JWHBp+aUu1SIkOXRhVVEEa2iaHCaYu3j5+OJzoD8d/bHe+KOLlK55pbMKwzUjXj3A4wt
rHoOE1Dr8oIoce7SwR/Ax1xkJT84n3kG2xapeClqekBbqFPQ9k1AMacXk3rKNzcgnrgsL9dnwXvD
tVI2gVWKUD9tgeCdt9f6rlraadBICvfL8l565oCstelXlHYpPyAwzTOxX2WFLRQZoc/M4le7KOvH
e0OxU59x8lr7/VSi7d09n/I2B4zxLa7ehXEo1uQ5hOEL4YP6uIHjhPENujXbu+8EYl93QrdUOt7x
AWVLbi9QFgabEnEKnlheiHRilrrg3k8COcrrt235TyqqY7sgIWmYWu7PLTe7YKSAF8ccoz16ZOWg
k3vhgb+GJrV+IAQRRtaFty+psSu/16WrR/zzIWB1JMjS88A+R7d7II8zvcAO2/z/xOxAOIURALnw
WqrwfcJM8rELsJHHzyD8l251NXsdn+O8NQMo+DrS15xWOVmJh/Ab06kot69lp71WJJ/0RHNpR0jP
74j9mJ7gFomOse3tAuJWAjWWrOFYeItU/PPdYAvrOCAeFW43InYgZfdQL1rDFIEAq/gESvFEKrO+
/09hPVQZ/DrbQBrj0jXk+F40fOjlqKUXZxj6mc3TqPJdzZMeaz5NMXAAzitYshniInm5GKXOQ6Hb
91gRBHhCj0mIT67nYlZzqShQE2STo0MXRKmHtV6wqfTEhU/hyml55Thx12PJSV+VTqugStyetBtH
+YdbfnuvHy/OW3CJPOUJOi7iiHh3lPkFuLOKPCT8ICYnUw2U/Dg3d4kSof4GJdO3rp/TbT79xKpq
lIkfWCZjKs/9d0iG0zLhBoCibEzFjFDVOAmWPDnsZDfQO3/1kA9VvRggQm6gCmvvEiu772JAFhYo
di7oeUJFcw0qOcgaXbONehyPplpUHGomlYgBfInvC0Xg3oNkJKkxmH6OaNx9gfKEbZ53lXJfzgkq
G7dcBjUXvDrgL9e9lAS1Tp0OarwW8ZCVhgvbsabSaWk7pCOuPt8qtG+LEGQrQp3GhjYNZn6yL9H/
0vyluyV1IQzD13BEC6BVZ/LUe8Weivm/Q9WT/qatg57gvHS7VJp7p8k9C2xYPWJXQgG2D/bJJX0O
WoPu44ficV8Pqhcb0cY1rElldgR7fHbmEsvK3dwTU8XGWxZYk4tSXaUBwlbyBxpzDJShoYZsx2Wf
XnFaENCrbKM27F+Mk95Bq9Vc3Uug4Ie561wgKjVouxilr96I2NfE1E/a1dECgpkJlFlor6i36cLq
XsbE2MyA4ywT3gCXqeLO422qOPxb9aMAaxkdtt7VmzZPZYDPm4VAfDUmwujjULID0IS46Tqaj8it
D9Zn//j/t2+2ujSnU9Xq7AKk3qPvctUbk8clyG4vynDU4ciS8NpNlISex9jTbwyM8JV1LKfPMxbF
FO+IlamlaHATg4N+ilWL8TDG1hdO38SLSSGBWprZLn7yzdv8nODsIVklWufqCb4TYwPqq4iury97
w0iDVdNNvXMB/XPSclJK+K5GCRZCm4ZfUrtJ6/lFPMo2EwSD33+PpIWOC6xktNoedrbqlV0EEJJw
twS1sDq/filME0RayWYdj81ybwlatt9w+0NwGvkqd4uzqDyfQfAJc3UTsM1a6hpbVDzI7rY3UUh9
QfRy+L1jup87GsNFAwzq6qnnDemPVht/vMCQpP4vo/kpXKnKcwuRe7Mn2QJor1ipk1YBW8cWOwpp
/KxD9x/igiBD4VeYKLe40RyzO6xcwfz9EZU8fbo3voKfpxNZuCthwJARg6nVeh9GWgMTlZUClyPj
/J5dnX+3A6Gs4NVpbDXeyto/0x0opwuUvhEtw8Jq54tbzIgcHAomn6ZIAP3ZsCYzyNlDfCGuXPFd
qtPAj97EfVf5HAUWWcMpU8lYoW4IkvfuypWBuaqbSnXwVQhEb/xJVTOptAxMB1AV1A/T59XJwr+n
hXAMoisDlIM0l9hFz9+k+8XtR9jdhI0xz0gCE+cPrLc7so2VTbFHa6bEU8BRKKQqRP01rr1mtwDW
pnhkyqo36R8AYmx8AhlpL0wLitfm9887wvEHN7jVJxNZlihhE9He/wKL6PvoBYX4yJFJ6M3MP7Iq
ujwRVIKDQ5SgG8LH8Q9eN75QzK2XpnRcbPw4X3BjIboXGBxtwN8wbGNVxuIJD57KBEUmqDzkmF10
VRKFVpz8SH7goDZvmLQB3z93sxV/1cCUOK3JEcI+jksYAXtuKuCoj5rNb6Vzs1iMN8WryLBNi8Om
Ral1b6ziHSrkoS4MZlV5kRxwSeYtgyiQz8FgHKUnjGZAWMfMf0YxuVjkQQ/8hFYlCQuFAr+qJQoJ
cLCtiYPRyYRAV9wjHz0Xsrn2Fn33QEdE641BxFJYNQ8H9Sb9IPcB3RVpq5fn7Wm3alABn0qJyvnJ
vXexNBe3rSNVZliVpyhYiGQTdJQNN6owRGyNBrMKKOqhysVtm7vbT2HUlQ+iPNx1HZdOvojiJOme
Wi+rvKulDHFO4Z3goEOzuVNj8vjuHR+zVxB97pN+iqFNL1Bee50Yl025zZWzbSFA1b7VETH/0lYI
mTgGlAkNgwsRT0xf7uqRg1uOCMCFEAtPuowfaZqCBjakCcvgwjaD6YcDdE3PaeiRzIhTy/bcF84b
bc39Xc9CH0ke7ImvXgW0RPbzc+k8XBZJsBoHRSc/ONofSNFhLayqs0rlI8NI97xJNtpSaFWbP1wU
kReiohA9wSShwERDdfPTLKSWG3i1JUXUKvNFC527xn3Py64qu2quv0VlyGb1hTGI8+wTLFuipD0H
xNnjI8DLph8ONt40qm/MkAwsOXqj/RrplzPT4PJ4RgXaiC2zFWU/XX3AtSAwPungue6ZGt9PKvBx
orQPq8DRC73E2jBV28NBZRuGigfZyWSrRsMsG4ixFLzMO+H4+z/ECYHfByrO8Hx55a/H735WbrVs
TPXSfV5GRzyGOEswXjU1Pedzt1vCpWJL5LDqYrhfBoJ1vKBrimmYzBhbG1rqrRSuS/v1RF9utfDK
BNr0tjTPBmW5hIUerSv/mAzRvJ4dHgVuFdc1GWdEBLzKGES3PJmnrmYy/YNjX7LUCMDFG/LCod29
n9b/tbHlunRuTPX/8Xg7tvFBBaCwJOKGJbuOjW/6DUjFg7+v8UkHlCZdupSHxaLF8ahW/TlQbt41
PYth182PgoDKbZ3ucydv2jzXumOyeOrEaylQdtwdcwoZAuJkhuKYjkTaRQAaKXcK04V4iub7Wp1w
3GmhpjdDmEeXBQ5WB8qtgEN5O3OGreuDzmzHgrgKrmWboxFNLjsP2aARCNeHNXFRfl5ntutS/XiC
uICHCssg/RzhELKy3/pZJ1iJ24WO4wy9/kF1SvliVajcLP2oSy+qihvQ5/nV2qiM/1y8I5yG83w8
GI37N5SD2/4+P2eew8+8nZxnqMGuSE1tu+D8Xe9Orc4C3zLorWvSV7WAhFxbwiPbu33KBo3858mL
XrteEzEIh84dC+m/lj1M+kxI45usqYGVKzlUfNfg6TkHlF3Wf8qiUC/eZG87xH9fh0Fjp4fOCwOY
XPGkPqC98CGJVlWsVLc6Yvxk5XeX4vnWy0DGe4d6JKZFv8vXD1Fc4UDQTRuTVAPPtHaozbRA3MIO
ChhdO+axqo2WkOlf5gViufXHToywrLRMwb2hmqHwGMS8b8tAxXK6lSfCdaCH2BUEz7vzDy47r1CL
my5nZ0yqAgtrfOWFyVL3jk1supBzViv4Cy6lkzV9GTxf9FqwVpdAFYvfaSEuIPByQJUCRtm6J+X8
u95wUL89/YDjd6boJHx9ktyTGLYaa/gGE9A7KZbB9FglCKpONKROW6ZHJ0zL0Z9muP/P9H7os5y/
oAfDp7x+oPwrObiSBJDKuxjmMbTQpFFuQ0OFPXsAwv5417FJ7KtNeJOQCRbYfXVKWgNJal7WcGq6
9w1pamUjj0ZqkPdZAN8RUZAJqWF7CpqxOTNp2noyACW/r86wo2dkNzmm8ClDVQIz3r6+VEKQOAC5
erDfaAISHO0aJbpAvfFl/OrXD1BEqtcUXGld4So/gWcXICH+/KXDIes9FPP5Bo4NpTF2EkSfURLH
ghV8GP0OJo3fzndXX1ylLG06shYV/i/e8CGgjKnKq2iUrr/NvV2+0gxMoEtdGNxZEeOrS2ldmkBG
zg2PaWKyE5riROrXAno9Xf6g3j/7UeY3SswDyVF3p77grQ9XTFrR24hepJyRrg13bx3wFPDRwNSI
SFwdOjjNG/WSLkRzTRbL4LJIURt1zzKzvZEwbZDcfm1IBYCaL1xveeqcJKpAkRwIDhRwLIUTueuh
KM95IgnZ+pgO/L4iCTer93fRcKwdl8x9p9VHA/13DE7kDHPAys29gSBaIeBQR5x4fMismnzBlJRf
IVoRXbq9vxs92osJaXCV1EZSOmG/FUgLSQXRZOU0SbldbQ05quoiCaRQXe6q9YHg7VqhFmFdl5/6
lV6FmZlSLmuq0eVgvCJfVH+aW6fEDToQncnctuuOvDR0r5RMbjOtS6PLyyWM6ImVLdOFBYndZmgY
4j5pulsrmer70GyffioyE4w5efrOkgt11DB1Z4tGpxWOXiAZujE/PBeU2YyOb9sFXs4/ao6tGGkv
e49/rn1g0YXr1BFYTP6DaFTFMvAcGus6xzJo0zKLoTNbAvrLEDDONGu+pHkvelxkgOqliTQFSH2t
eUkDcTGrLS9mPHOwfySDhBDEIEg/xLJ2FAJdW30rEzp4Yw5Q6Y0x3wvigKY2f9VL9UxzGfVEBNPw
RUJjktojCr0boYFJwfIWcSMf3JhxSP2wvbOWu9IHOTC+Loro2651/W3JmIi/jO8nTIwxcfA0eqgz
bds3D6qNwRAF77FBZqAhPKP+tUyTV+C4BBaCpfsXnw31jYPJ8arue7wpA+pL4i7ns5icjQMVqLl1
ZxWQ0Iju8HkfSZub9YVttX5nEpB6IMyK9rcSuQUHe1cvShGMCGpIeYnXviOWKLtfnEW8BgHMTcMW
DViNSo8x/zrXEsrYTqczdTMNOFHpL/V/TpUSDs6LQliV0Phgxe7Qz4I28WmfeGe63eW3A3VDo1kA
jZ9nSEKi6vjT+oqAOvH1dKFUrgKVt3FjQ1QLAeDPAH2vGtk6CCz38r0mWc5ZNf7D+drM7g45PaKt
sZ2QnZo9kSVGgPXTfToZft5oqgQ9rpo5AFa9t70juF9sgBpuvhMkSqrlKRpGJwI9DHIhLL2+EODN
0WQ5CCssGp2+2vIXVuxC7BQiCIjSpCpCI5ysmca5Ul8NtlAgkeVSepmEyDQPIR/tELopCaVjM9k2
Qp6N6tZjKW4DR4NSX0Qjd5qoQoDhlT5ygpy7Jb4b1IdFJHhFV0eObP1dDIzRlCxoTOZ6dzNuknfx
51nqtYw/xu6B6faZ4zoLIMO9zlRNwTPGv50monfCtdyDs8KAR4qB+sI4iU2LCMuq1/whJ9+Fo317
aUirfTSI92JG/KqpGNE6SjpotEQk539kvUmgxyV34JVJOJ4h8FEpIpoHmNf6lhccUxwQDbMvrKbn
5tWsKrhaJQk4ssIfLpcmHQkgVjrfymhujxqOQyVWD/Pbo1jnpk7uD7VFTnmdOkHUiQhG2L4hg0J4
6xwZW8M+3oZmavGu0g/ob+69U9zdH4Ks16rDbHy9wU9xWHuxdNart02eS3/htRp+6uUMqm5FLqD/
CgNskagRYCvt7M2mJZLVfiUwUTGvXm/f0HBCR50JqLUckJnCbQnWYhN1dl7HhE4WZtrkPv2MAxYU
JlqdMeR+EqpR+Q3nWFXHdfDpOSL+Q7G7rTUQID7k0eeTaU9m03GNDGIkLxik8k/TIktjkIIbuQjQ
Dk+0HWXBoIAT2Xyo04lXSwJKczKJhKrAFhNDEQtba62QKoWdtfosi1HNgTZitF4ZQHTa25H2XHoY
r0E/t/4XkFFBfE0RlKhaiW7jbrxm9LBzU07l8tRcyA8OYbKNsJ9ekRfaAj6JM6NW5wpYcgAoCpAD
IrZafUFxxNH4R3AXvx9c8RzPITxvDoGFtwt8EMlElXwnUbJLV1rpHhfPC+OkcGCkqZoDl+nLOpSF
MtDRk7vlTU+r+B/QkE05eYjaPt6TnbvW7gM4Kwbg6ziP+8yVrcipDYJbqkmcmbmF7eRjdgLZINgm
m0S+/7kqBAr/OkyhRSkcAucT5Sdcvsl5qLUQyP3b7CBUvsIHfXozaYhBkE3ec7PntSCGnmSQ+vTC
ltKLQYujmZT0Wu84wx1W6wCjHiMy1rJxwXLDuh9q78QFGgleQJMVJrVxwdXjH1YVot2ogu7gkpCg
nM2bm4RBAywe2vhWA3ie5wW3EBaZAjM9rme8EDtSJCMYvZYyOwwOVnwOhvWo1Xkf8y35qu/tefPG
sp1qKQFlicVBwymXfk8BGM6xyZLU3EGvvSnA6XVvQ01iLjlvL8R/fILpoAXqOc6PHKDkwAlO4JIj
xL0SjFDHyeH5TQNnAp3+M3o+KvRc0EBN9pgb80JOcjnWLLW8SjVaV8P3v8zJKwVy+tTlTL+DDQhJ
5S7wX2+jOVejOVGcezyRxlxevOEuzI/mg+y1ihQxk/FMHyAIkXAU+xI5B2xbPIxQ9F6C2ccFTffP
76T8dIdn2zASFAyZaYmKyp2OTc3krzBs43dZwu9dgk7tml60vsXi3fO6GtdD4ZA9fh6SiCWVqYYp
79DcAGVVACwrUToVsWXnusSay+LT7SkXvawWGM/v8bEkP8o1Q7EvFN416bWPMbDJNPUlJ6uoQQEF
PGNnCz9ehrpfLJBm4UcYcMv7Af0xvpXM4DYaQ6m6XFn0cJZJfIX3gB3hq6hgy2aiSwdJhTZ9OzQJ
87GUYlULFj7garsqvkICB1VWmDEMg25CdMJM3aR3XSo3tJMC3b5DBaubpWVoIziISwil0DwMT3qV
dIlA86hiz9siSrvTaG3SwjRxuqaVhaLJAv4RbGh+dBuH2dCYGQpwikYBg5Wr+hotHLTV+GcADMHD
v3lH7PhP255fYpvAfVlbYMrJnuRJaUyTOgDJJxJyO+xMVwAuOkNn8MwobMM0bBFAdfAX+jY12guW
2hh0vDWgmcViPa4448ORCfYt10KgDB90RylmM6ClVHUX10NHkzXhJWCrvKvqupgIi+/IrryyRIw/
PmVaf0B4Ys/qEfLdrNRVxteh4ypElfJtenA16GECWNXPeWsvRZCw/wZ+CAAN04uAJMp1zrqPbk3W
mwJl72WpBr8LmaQgXXDXmqVxRyIZ/uz2pK6Qn4mITvyKSerUGSQV0xBYIxZ0llyeLMur3/2htKLt
e89E79pWEQtXs1yiulxUAuzpqy6BNmAlitCFnhWNEK0bXk5VxNu09XOFR0WcwQ5NMrrjx6N0x7ml
v29NwiyWWDLftyVb3MnKjZMG5KYEjUq2FPvjQZDpRjoKW2LHtDV5LWii1KvrL4TFcoQreVf1IocM
SCqQVE+u9tKsa/S4Z7irHAnA0BcndmT7fEAXIvdkrOZkVQvmjGexb9HmDTrNiCm87ixdRW7VT72y
CpwEUpm2oCnos7HJluTmRYk797RgfAEZEn6+bx4YpZam6DVsJiaPn3TnpVVnwKCYSzKbk//INiL1
LzIK/JLljrWJyl1fFjLS0Q5qZbPfNLfEJGQumUzaIqGv2880g3AnyaqbowZH0Az9Kvm6FpFWvxbY
kZx1fJSnU7xpDuX5jE+F2uW5BKTmf614JaVB4Ya2LIzFXmuLsBVIzhDgV959HL2Ej4a6dw+yFNo4
nDpR80WzfvxrJIPErfg6hetaX4IjyNZ3G+vTGNOayTNWZcqI2q5Bqt5UoNPUOkpFEeRSFHydE8vM
WRrpk8ZXHW3nZIxbUebhym3BbLEV0gWDTQVRFzCEgm0YJm4pjNdsRpBTl3/Nfgl/wIvTv3+FOi0+
rzk4WY4MMjnO8uSxUhK8VNCbsrThboKXmuSom17i1mHH13zftXO2IMv68ifaFHt45S9Vmt6jR7yV
w8Vu30dGxiM5K+OfJSmKdIPCZ1bc8Slm9UpIT4TMaIzYnaewhUq3nynHMdkvBbyzNJqUIgHu2DKc
jUEtn5gIQr7DmT2ayWz32A9povm5vS0bVccYFZcZomQQSowqJ07De7QGbNK0eWQUrMkjxz0HwVeA
FRH/yYPKCl7lm7z+zOKaVdEHiezUbgr746USrgpqMZ8vaFrYcudFK1PUmQ2/PgpGm9Ue+p6pOLRW
YvZ1nGuOgOyl80ZSy+IZKhnV8FsHZjLJtlqrdSVElB9M1CgrJrrwsffxQZwtcLEgeNuS1LZieJyM
DdcbJRm1BYUW4D47KGl+4E6/2IFbjEL9ct2yP+T2TFgOfbqi9Il8pLZqXkF9ueezUUEHelg83IXO
J5E6dSemDHgijxnRelEc3AKi3iH8YPoeLlRkVPF6z9PCqav3BD5Kq5BrL4A1oZKMHgBY93NKyovw
ds6RijAMb4IM0lKgWfSasTLhTgpNBIOAKLA6qWIdAyTh+2j0zTQF/gT65cYGAeFgEke3va6gcqQ3
TNDgTT0EKNqByt2flthhgZDkK32Gjc9MYC+cT/uebGLSxZ0L+QydSv7/hnMT4SzZa9o3Lk4Cd02z
Vm9bjR/BaZSFXZWLVigy2KvzcASHPjbmWRfKBs04gTC3dMwVoPi4A/2Q3H3yMD65abvopG2DzJmJ
yXjZ36rFrrH10AsVUSvvpjTJwOgN2qxsC1ACnDkuYDwv2+mqlKwvwwFMinj0Q0MEi6SEqWlKySSl
+dmXl33gtJ9HNDlbos0Yvy5rumdbypSTSFHGZOQ7e0fkpN3DK5XGrGqWjLYAli8fQZXhngdRHHzi
fGuKjW4N6Pi5vwgh8ybfxBEaKL81xC5WNhvR4uT1FiDf4L5HccFA79ck47a8YE76PNmk/0XXKTUi
cRkJkBJdw1D4pucjAKcbspt6T2EJtm32HaBEFa8Z5w53yyDzvlTJmnt/D95APqFunb9gpz3PFFs+
8lw3yVzt3Fc4Z3Q81SZ+FmjV6PfBctPWKkaQYSljYTMiari1n1KFWVfUZXoaibqVs4KAwWshCJRi
aGDd6m6/N80yFACNqd5YcWCKwYvkAQLtv5pnbR+M7BnMhOQafiCuPu5tPbN410604i+WpkFJ5YHE
u43WXnz1RWJr5ryYxmmqQOKjE5cz1jPHLPl9XIvHMV1Hv8JK7K3Dq6S6EBhv8zZJimQ4nh8kULKc
/R5Y1VnF/BdbnqHgrcD+q4KbjqJNN3DfDIsGVbdg+AS4G/YKh3Rz8Gcol9tYmVFQSdRoRFgm749Q
tQGxX0vTkO8BF070ZWoK7CdKtche/PLySCM0luy1WrxlnARN2HduH4/N+ltq29JeNsrfOwROiJ7P
SEryd1/m9ZuDUn1Q0G04aKLeWK+meD991d6Vp7+IV8TREi+tLT+3H+9a5Z3grn8cXmrUW/wavh5f
LCxu/qRBb+hqZ15UBdRreBE9ZZoJtSjzMTVf0hecFkHey5r7AhPwW++21DCJgq1SvIw871vLVWBp
/ipamu3HN/Nl+JWduiMJwjj4OGY9un9Td3j+ky5jDSJR5ZfRK+r8A5yQchvGKmVWEXmqQ2DfUjrY
0l2oBVOMzs3t7NsMpUbP3W9wWtXfRVUwpbZJvlyKAw9WdZDqsbVOblYboGnELeiBTNzs9wzD1kai
czbGvQ205UiDt7VFO58xlNfIqRylmVarvfUawzCsIR2WzKTAIziBQlXo8whmUuMrvKR5p+SiP+I4
Qk0heoMOQPvSEMslZ152dytdJKGVXTIEY3nek/7puDoV7CStglxrDgDCn1n9GgVSSZcBdme6/rZ9
e3KNqr5YfZuZ2bUCyl9HVA5i0SENHI5xM/WclvNeGXLparUfd/9IPnoXiOrwfPYlKRZPPNsXr20Q
uEQnYcUHTENG4vj8rcyygGqlvLiH6F8tEesUr2N8Qs8H20EQqF3q/v7Sg3fkVbvt7UUUQrHwMNzm
q83JL5xFKj9E19NkWqyl7D6cmu49nnquJdOY/lvFKUOVFK/IK9zFJo1rovy3SrThbTvlSS9Sn/sU
QvY44mZfnlCeBVkB+fNFRKV+gl+3jBJJEmH1CkwC2YNk4QjohjW9hDVxmf3U0UKOLLiIT/Ma++7r
Fy5Q5GqIp+9vbZGpAvDfjGuDJLFZ1WgRIzDrs+hT0KrqwZ3Fo83xthzum4l7bKtZq1P31SRhd4UI
qHCHEuNc/f/NpW2Py+L2lHXSj2cJ91mfPWH9Yt4GZBAfq/wP+W8s0gWRXbEmKxGTY6iW1XGqvNLE
sU/VukR0NAtHY+CNWiXKa98+UI5P2+nU72RhbgeeIRgOUlbrkK6YzKMlsuhpGnOIo/CWeOkXCfgb
/bDdC7s1VMAWzs4/UfyE8F9uVSj7XkAH70TlwKfLiU1URtkCnZUg4k7qGel5KfcV9q/BFNoNEyDe
3RhJYms543FfH4N4ANNjslZ1RVODaKu9pxeVQkjo1wE1ezESr2QNbjg2pQDC8WXWtTiZLm7kz5Zl
MTcxkKRYEK4qL3er7wpFYmqTQpLZ9XsQt8OnT96+JgvZxVGSywOfLLVGljLZCf0VoJpr6iBgefz/
ijq6UloO7rVdsfHWTTFLIXcdpFqZ2WBjWMgcnyt+lE1Ao52wHk8dDzFjaF4dcAGX0XkROgURLiIy
8M4C44O7YtRK/akR6Kpbn/l9H9mbPOEOM9/iKgO7y6UqYFE/alTGx8FAxH2MaqH2LZS3pdds38Zu
PM1azV1WswkuZpMorU25DoprbtHbwEWH1hDi/zjiDWkaHCRAMn3n3mmUmrLmT0NhHyoRVOdkOqOD
BEHlX32Bnbpkx7oqVO+Qw0RkvKzGMx04lYevBLe2vGdgeFEEJQdfrwQHzQlWShrBreKMDD+R/ip5
s0Yes1Wjj3RO9vvXcWZZYaqaGsuWLJIS06s64/92BbfVnJ1UR2mVYkrSxNCXRgQg1kTGIwPC+3WL
Kq4wCtc89qHQwm63GVDbj6fg9cmZAnA7D2uOne8ZITPqfI4fXh0GtpUnDP0zjuvN5NvFiau1f30q
O/4IE4bwbq3bcZxZYc+wnkl6WGzUN4HT+vrHDiLYk9VIyKOTR8+jsildSq9rIGmnlxGKO2Q1vA/8
tDYWyuumABAycaQVOjfmp4/102gBk6iPTCZlJaNak6/xb9ibjgJPPfCHGFLEOAA6byCHITlFeD1p
DX9Yl2vxBLpKxtKSP/KyTNEjWScZc9cgJ260IrEAL/0yznCtSwishxz2f7rIMU6P/4G4esMWXXQZ
95KdU0aPy3OHjo9/wuHm+sRKt+FVpnk0Gdid7aFBo/xIDudWF2Lc5XCG/sxPF3QnzkRYKNg/pjP/
U6biSaJQ3D1QPLM4J+NhPYI4Vhy5Nr9nS7KbfW1v0QVdT84TELvm/K61kaseySXR2mpSj9LzTLxG
iUOCrE/k76ikgCh3vkzw+Yrx+irf7wn8omSTiLNDnPNkjSdgUeoguvNhsWMAqSxEx/6x+MX1OONa
aUrU1kaN8Mm69omz/t08uhq2nYjBLv8a6Pe0TQeJx4KQPzRjuwnvygRi7mEvOmLdEmOkrM/72JjL
9NKZvadjfIREwU8T0JS3thEpnUgWeGHVd3PeXEtm+cz2wtZlVKRFwPqcVNPmlF2cb39j2bubLRco
GyfvnYIylDIxI8LhlZRFJ6GfShZ5TwuW/nWCYwrf0V5h/L0PBm4K6p7b/XqSDNMVKeeMjahAbpfO
A5wQW7mEfZrKqiVFz9R0wmBP3XKX+qRQbxVRvvTilIY61qAZfoBaCgAqizdyHcIHzdeIbLhS+g9s
6KD/NOBeEuiOoXFsJ1mKLIefKFMTiBz+nuCLvIjhy0RZkZDQDjkss8OOsSeak9B8NC21rBgqve7b
Ui2AYZMfRU3de53l6IBpIKhtNsDnrcEgVT//0p4JsT+ZLdrdaCa77y8M01eyM5S12+jBDyin0TaT
LVyxuZIludXS3qmL7NywY7dFeZVM9Y3pYSUaadhWrG0ssJiYDrnitVJ9g2yVz1YomVe6UQctJJW7
T7C9Pn9uLls3iLUPuZxFR3/1nXV96H84KZHVuY16UbTCQLMB8rtjKlpmc/g2yAoBNv7CHe+SpDBl
JE/MJWAg1XlLwSg1LbruKN64ACY/b6w0jSdE5wEY1AaVmx1vNY0586LOfD5KEOGxc996FMnsvuKH
UR0QwWkmsF90i3GDIHBeJWChIq94SEPeuPO1ZcNrTsWIjR2v3ZRFnZ301XGAalUOGmLIHmQmXdwh
3hF67a45jiua5HgiV1Pd93wMwbfsKZqBniaanQIxVBQHW+BXzpVy+WK6scnc0zfLwx21G2QPBha6
oP+bcMFQABj6LliDJTEBIWWdED2oynX/gU4ma2iMvLpEoxq+0t6PFZ94JHS34hw2XHdWVY2jHOil
AymsHdfOgrWqm/p7Pij9r77tYSPPTvl4FSE1QxbEVu0Etw8trceBDbVa1239aVx9Z3J7SHaouVkc
EFePSrqYfnMsX69gpk/22q8cWFxJReoUjmy6GCtzWQ4q8wUXzAcknKnrPByjh7TxKUxs5/2Q0THr
jphQjFHCKyPiy9HQ5RDVlQyq8dzeJmzgmKZA2uctiO3a2GAzLY/P3Yvl0fEMvI4KLUQv5uhBIAXC
hZsNWz7RVQultASnkMeh+WNdPYzOfD2x0w6IliZJ+ZuANDBPTZOcYskq1nc5RDvekv7HI5++DibL
huRXCT+O5/qGU/pDsNwDE6zL0IbZxv6Mhlzpqyo2nDx4c5Ih7ve8YysfE745vLMZtCaZSFzEWJZd
YBZthb2T3v+gb4Gqn6AO/xt4M5+wjMlO6Fq9UmXS1ZURvPn2T4WSZVZe/prZgZCY9H3Q1GjFyaff
+4BPuTJf5i96EainpRM8e7nYm+SihD9FlK3Cerh3er3I6ezedDOX9j/vgfUXQWXOYzzVGk3p0JnC
L3RUNuaLYHwCSuSBOKVND8dS/u9oKU5C0xJCrzuRtBrh558tjoh9wbZLil3ull+BmoKCAjuhdTwm
HLVdUReemCZpSlV1Dhm7yOYPXaJ2hxAWEPTbE0eraaF1TrbyQ06/k9IpGT86iqxuarX5jFe+kAMD
2TW+pMuHW3qA0fwSZevcfcVv/i8ielqTPMIx65ju1tiTXXPFFU5CXD7Sdypl3n/orlpopQplpIs4
HyOiDihmdT9RPKzmU13IYk91D0RWoI+PyUJZNwvthX6ddClckDh1T0bC7D9KS3ekER1Y8hOUVyfj
nBiFD/LJe3pa7M525vsUGSuX+Pn0IViQHLw0dveCOB5gsaeolXHxYXgDgubzFLIliBtUW4AwZ6WF
g2u3dJSODlwiSJ9eKZDJBNBCtJ6cr2av3YoWdC8YQ+uAvIXJlgs+vwHnqW3BosFwmWSG6vnOH+8X
EDRoRRmddfv0YvbZWqSv5+VpjASZACfnPKCOJRzcKz2RePRkLX2ZeDU6AhcbQpUJ2Ur93C2y0X2R
veQR6WMovo8LQ7Z4ydp3+ERvBJlNro7KCzRn33L5QPQo+Wlim8AoVXC7WWKo+yde36BeEfzEtkrW
PkOxSwsdLOPbBgUb61/wNbEGbUTJ7jslkfdHjta0dyAMqbBh40BEx9hoH1HuUp2lXjLNwnLxcQnJ
uOxGrqz9kl0sq09ouL9MR/DzwuKoaJcTehzkTAdkJ1nFWKIy66K67RnmvKsvdzx8IZZpCW0qUcBc
AuI3citsaqav1xTBL9n1chioBqgROoLnP5lLyei0tIfI3lx+zwcpfjWb3xTVztLsqhkUkwehimw2
8ToI51+ot2vdIKre/O7gHTi4QT7LfvgugfzhtLIg0kahLwUdTRDYL2jHAiYRnIBc5OTT5bmg2Uwf
mBiu784TpyTDsnWhZck7xLm7r+yRdCk5osJajYxokENT3GT+4ks6n1ISC4ViEYx6tUFUZVsT+8bF
gdvN5LI/oWtS2bpfwIZKN0HaTbddVID3fyPjMjg3UZHCwiYs90JXmGmZhnZw/QqDn1HSUMz6WHag
zSienwj6/PljwtA4E9twCO/Jd+ZEWToG8O4DXko+xWnyjc1vhasGC1nQIo3jM9Mvcf64Ezoz/2dt
08qhhRGaYBpEX8hdY3hvuDdHrTjGP5RdTApkzB9PKFPuYL1APIOk/6FSQ9/P07yco2obiQpTDDFk
9tXqUq9UoN2JqKkxGuK9lbH5KM/cOA2rtZM+OVzbB+DG+aIvvpu76kC0ggg0OKE2xUtiqjfkl2vd
e+lHY23TqBG6ba2l2Uth2gE/u09iovJbVrem0r8HtiXTBoQi5Ht9hLKWXYV+7fC0+ix3om4/A1pU
JAznQ54pJVhsl2DEUrfg5bbkLqCsnw5htSzIilflz8usndYaidgmAQ8wQL8zUlVP+VXVqvUpMoux
THD+O8uUoaAKnyHQuWWv6nSHMJRSagPLEqFzp+xnhXDtx1OzNwroIJphpuWiaO5vCHt7evcoi0xb
az8NxQBxs/YeVClQg2SNXM0vqi8Ln5mhN/QNxnoObp6REFFDfo9nEnWJ7EBvhTrlHE/oslFrings
Fo85V+LM7rhr1jahN6xZq6wz7AbLGrOkz2oWRAmyhMTHpQQa7FhbbYJlL9CHyDD9siSJwL036RJ8
dIRxyD8fJ+8B+0Jsx5j28WAoSdytgdyDg3ecTtrs18GvYGXXtDAqV73/aKFezIRNAdnpveanmFUS
WC54GK6Zxbx+F/wZs4Dmzmhnd8IULXY/24qHfybSUzpZbEPZKtzsZO0sxCGhil43RvEtZ8KyeNWO
6KpduJy/emsqBJ9jCdQndKDePVlr4wp56bQY2K18WLerNGEoznLEFkh1FY1pwo25JTW76U8ZFyde
E0JJRjP6ZupjFm/1tdI0KT2F1eYTszAPTc2U9NWPNqxpzPgD+nqZ2cdCGtloIMvE7z4wz9ptq/xc
CRnPkBRyCBBAQ1ycHEJkcxJF9goqCpvAPMf/Aog1ozCixejfPh3G3OSF/vYcQMs4ZUpYTdpsALNS
9fGaVO+OOSerCHkww4ZMkT9EpgzFBtgdLg9fu+5Ujuwe74KDiMGMrds8YBtl8S3hvdmf2KNAd1Bw
UwV6I6YgZtoIZXcKP+LAsX6+B3fKUiPrwwDuKnedOAnQMQw5k2ck3lRUGBgP9xZzWWmRAUixzbA8
awpVraCMVWRzy8KiCbsZJqd6hO5UD4gwUFI4CzOoDRNgpO7tlo7sfdbUsz/KD1/X1gb+nroWP1EC
8TiwQ5WoitFL/x6iBih8IwWjl2xLSTAW4RBasAOKEzS6Q3AqWAaSXofj7skBLyBjLPdxZlj5MmiA
YUabq+hrfVumsrclHcAGBMOoLHfEnrB9X/JsXALKH+Zw7CGqq4N0vQ2X/uqpcnQIJjaubcdFTup5
h0+QrLDoR1V1H6iayFQ3AI0K76doIORjORqdTxjiCDzgnNKLGsfHvGx/6aT7154hz0XY3wbk4s7f
LTAw0m2J1Mz/m7xd8TGK0msXOvmJuDdu0BZyxrH97HmNAU1CdURcrGx/CY8G3rgHmOTj5melcXoU
tLtXAbekRTewJxiltg8Dzsc9yttjczNandE2kki5aGRE9yTf0JPA8YfaQ5UxjGhB9I/tWtAobEgm
rzV/gDVz8lHKJEjfWKW9Km2PbUIA0gxzZOgbLlH5zMctvm+1RzN0xUOBTIvEauaxAdFgviZpy2kn
TV8ZESjFYM9g5ik7A1sVxeU5QCZqIuJHDG5lth711vmJCXgYtlJE6LDsJfHdo7xlb7eC5sMwJPdo
dg4XmH3HS1fh8JgPrcVcobif+tvzpZZ4BDFYDN1GH+9nDEvrI65KmwPX6UPVGoYnUO3yP2ed2IHY
22OHW937JN+WVN/kE2JIBoIrjBzsZ2OU00lXNw/Uooll/FbiMbIhtrS4VjYb6TrwcADLeUv7eRmc
URIKLr3dHSOl1MhVMGxbiqQ7yRqh/xwoPjcECIB+Tj1RzyGy/7yTfvjJUfi+BxvWSruHHgA24rnT
3Fw72SZMrDVmnLuge+z0lPy01pw4HV/ezllL9XkEScgHU+2mqAVud16BXDtEa0FVNIvRmwkmw/7m
6AOee75Q6XOJCLQP2wbw3JYCECPYMlueQuPsrOEovlr3jzTIy7s89o4IDi7NhaOPhlZJPUn4uBnL
WV/2FtmJYLMVXK+elhq/KnRGN4RHTasQlMeiD264P2nfi/uZjz9x8uo+aUcvhi3h5IBwFiwvwKEs
6UcBkQ/75witXa4MpmMWWDLjESyXxFz1JU6qkwB7psUgcHehdxoZh4RRkOxEtzDOsed0t/mRmnCC
KEV4j9Wvxk6gxpAVF9qYlQHLFKLp2G0al8ZGuv6buz2CQADAizMmS4Z4abqA0fIdg6bEalNBFwvf
SkMHtMOL8iG5QcmEhdqpshuVBiP4+IzKDECVVImuganTFN/wRP7syCTPal8GtMHYDSwUsq9tqCSD
9SJF2zB4jNkZwtjaGBQbz0DU9hhJz15JdbUNpT9pbdIAR83lYTFp8ZhNiMpFcSByDX5E4AnF4Gav
ZMjHsLUF+9/1NT7twPKCkPebya4a66nM2JJsHAelUhwrhTwHSJ7Rrtt5WIpcNbBQcJMSw2Cm9n/k
Xyu+duiTU0LjkLCkgRfczk/HYrBRHqU3zyYGYip55vjOxc6wBeIGlEgosSfJyLf7dcPvnRTiqLda
64HXNCV5KsrFPYzAy77t1u6dJfKTcy1SGo4wlC5hgjTaNlmVVqO24VK7ubQ76N/tabrh0HFE0aOT
7NlTmR++JEnH+TNcvfJehiQqzEK41LzXwSEdHIZaTcHIYmMDVxSLZjWClCPUlj72PxG6Se7pMNuJ
r4kzwQYi1vM0FQuIlYLyx1Psq4Xsd2Id76/sI4eU9bnvBCm2tWuQcnJ1825kYdwPeDVsa/rWzLwy
XBdQiNq0ingBBSQrCcgXDD2kXTieUNnz+kImzkOIltwkCIQnVwFHZPL57sqX01/Xf/ortb4Kvo6d
xKwKzGVfCQQ2L56FFAOCOj2wuqthhzX7/QlnEvNxjGcjTgZ3xOZ69hDvEWrSWZjSE1JmMwPQVOWX
dnuQXsGDjtO95clGF3PqgVLDBVq46PIBmOS9ly/kvCKuD2ubmcVOZhD4xKWsdFYhR3LDW8IzaRTw
zb27mDGYm64vLG3ru3CcbzobPy5vUI59ywnUWFXG3g7YjMGDz9mTMW1vfEmHvqqSytn4mykbUYDZ
OTJ8gUqN+KWKN4//IF2yCtDAVnJerVJY1PwqsJom4mXkIACLf8QwDYVMYFrwmH38QucIRl8y1oYK
E2OyPOlvsPrEhofs2ejgm5KabEQbEMiDaikzE7jqBha9yWRttr9cnUtK3tXVFJMU1gXaMu5f3KgF
TY82WZiOaOxGE/3zj+ZMTNe6+zCUO4D4AiJGQDKqME0rRLrXL5IL2EYcFAzlTGztXKZYkQto79JM
zMuNxXXS0yybAUGvqEgIO4OLB3y4gQzzXrn9F6igFRafQn/ckI+ILv0uR6jbF2MiP0tGw9QgIZlp
740/aifWT8ZB3usYjI2MEyLaJGX7vFhRTbmgiL5yXa35P049AoWECN8rwvwuSBB5l6g+a84goNsM
eudbgstPv3K0lTRl7Y5cjK8LeBzxcsCxYj71g+cquzjLvEUqxm2ElY8XNeLiUMmFmMJoD8IYaCXG
ZfQ6tkKyVuXitxV7Hp6041X5p9CHK7JOqfRfGFug0F5AYnDfxDe/RHGWkJk7pI1pIRd5m4CASwJK
5V0ape5yCawHOxzU4xJXBmw+ARN3lhp7PC+jhHlxkjCIWeFn46Gvlik7F5q1rTNaKMzAj2tsNZ5r
oKnvndsPCFsgLAxRjktJkuNSVUpnPBffS03KHdEDQ5nsRtULLN2qEHxkHP4XYeAyY/1U9jzQ3+nY
/Q1Z51UNkTx2thgZFndLIYzc4oMgtOleROKJ5/zZooJrrEFnD+F9M6fsY+tdpOAP6yGWcaIh440x
x3rP5tRYD8rjsJcireDM8PwbqakZZdNfobuXiW0dGw5Ox9ASTtVeZOcgteKNo7eNG2pMduSCfLE4
Ljx80hr0RMOCkwhF6lH+JdsREBtIayea7ui7WSjWrHUxGyaqAwr6JQiYuj7VSeTmuNT6my0lfq1f
8cB2vDCuZ3j5vv0w/ZTH5YLSOC9hnuDWymTg218XbUBwXynqdaGc0JYaHUUnTOdAZO3wINadry+i
fr6t/jzKWb7i2oI/SOYMnZU66v69NBvZkjKamLHNhTBgy0v3/eHlP9YuuPbbiIdFC3joandAxYd9
sjl+4dau/6VUl/RPgzkDmtd9GSF7d2EPKIakFOJur2oMdO9trk4oxNbOP4SFGbY2WT4BRNgDOf+g
/sAGoh1WPigrDiMhZYamxF1U6SjFhWo0BMgqPdJ4bgUpn60N/xxgKDtfiuWGBMx0FZEE2XtsRfGJ
E95GrEWTYSrQjzQj4GUEydCECrXAss0b6fai3KthEtpAD2Rn7Jw4nNnslusRZANrFvszvd4Tx2hi
a4jBnvLtyzC7QM410YNyadF+TUQCHqo/wc+9jhLQ6L6D4dNFK9BWZg8x8+ogoxSsUmrSM686MEaw
Cd1A+zqb+BMvynqtABKlKHWQnhcUTuIFM05H0UTURj8kyeDJ6/OTJzMTnPTm+02Lf4Hysn2Xi7Kg
PhTkowg7isaGOml2Y+IS9U2YESNeizYTRB+RZRb+T7HbTif1WnBn9XKsQWrvwVWB+xF8dWNAoILI
mRxfquQf/kB0bMHiw5q5AJZJpfrf6CWHHAbyjP5+Lcu/ztauxhNcHn6qmIWVKF76th14zoPHFSuq
u+y0wB5BI8LhqeWuCVMLEV19zUNjwnkevir/Kk1Zn6ijsH+ZmBVkY725bAQbWV/uHo/64rx3Ge65
oWmPGDquTBAz3lQaRtfLS4p1sCaiW4gqh9iGHqoGkpMMrUH57/UHzYDFdQ1ljtvZhsXEz9QJxUJm
Ddzsr9V71hCGPFiGs+f9JAPVIe3ChuO6yWlq0YLukV49L5TlbNSmxkuyyZXzYXXeL++AsUg5/AgE
1xux17N4BbPe2DzPGAtcHRNxYwd1Rk/ttqm4Arua7bi99/oVizNaDHAoM82SlSRT0gDzV70+InRT
Z991XjkIvSM7nIOcEAHYMoys6VtHHfIL7u02Bu7A1hHoCVTRCTaedq4t5mfkQOkW4XFQgWmGCE4w
1ces7ejvoC1fERUZe93UG6e4bM47uniGk+4Cti1bLiM8OKtR8bWawqqqP+9SCkUmB7GFu4sQL4Qo
T2y+Npoy6V2Kb0kaCTA9cIY/PFLOQYTLWHaBGY/hEMvOFodd71r6A9iBEup4tmt8SDCgkiRBoMZv
3IZFBtEmkSALw84p62V2002k6ZfLoenOoUMSc75VthTYXq8zYTqHxfP/976yWxoFs8XpMYiNKcqh
glc8wbz5yn0Cw2pZ/f5InkU0YDfOKarJkCQROgUbPm1kiPEFskiKheK9unwGjT4k+p4zCvPD7S+M
t1oi3dKQjDrdB/0MXR+kJF9dmbJSuaBclzyqzvKzKyd+RMIHOPXX6Aip7MNjr62+BONeSBeZPFCI
Rs90L4GC29Vw4in1rGWez/gAqlklu5Yb9l6NFHeK0DJO4N9/OP5p8AX+7FQo9dNY3pds7QTV4Ua4
e0iYFHwpQHDdS+6mO6kixkzP6Y6XHQJxGAzYnJ1nEq/nrIdHVjzndaC3oe03+5zl7X2rmeu5ip5M
HdAh5+DYREl6QJfPbbepY/6WpzvW9kV4j1KGVpOegPcscqmb0RIuRraa0UyN2vhDu0vpXW4Iq7jP
i5md2JXJeDvFpqL+KTnTLB4xcrWB0eDQMCERQqWWvSHq8jWOC7bxVx+KjSbzH+N6FOuAMrKkCQ2q
eg0xNZdanENx2oDb0hlkrFPMeUztQW14gyW8JD5zxna9wugIB8TmsPL0Xavjy63/PHjNPZM6M8Mq
PY03sqFTcfGl/XrEvX2UXbM50hLvP6NhiG7OK9E86SSOJ62RMweRc+Vm6DSC3mL1vYMEkiZyN6Yt
ZgdK6CBk1OwQMefo1Aczgd2vHlsWBSqDMVX8KpIQZwXMWuO2KvoZ52VoalHMF0S1jqxtqK2gjrhY
CdZw7EMQOCFPd0G7xqXUKMlTvH7ZW/4+ta/vXvk1V4MLOTjATSwFVRfxNjAj+zPs5h1ljczBswbQ
BAO2ytcwKkzfGwwl/slBXlhN8jefymQXpBJc90w36M10IIyFwrrb8qN+AFlIMqNy1s7/LPCbPhRu
3N179VxXhBKJj6W/HkJnRQDspffvgb3vLcS9nnyB/7IfTg5r1MvRuWITSJhTW17R+Q9M1L69wbW3
5pPhtm7Yi5/ehP2AT36yRapmirLsdW6k56URtby6NzGaWpyooEIQ8QmxZTogq+rzNgNWp+MIRZfD
V61cmmRcO11p36KJ2osXQ/Iv9s23A3oIObwgRPmi7ThyWOJPbLBgjnuwsGnPoxvjGdZa4H87gOiL
ckOikTsUP6Y/Bebyg+OubiRiIvmDhwSmDAUvZAGvzASKZ90bnh3iZZ3mvUkRlmYiarzue0cKKitS
KRD+p4yv1zO+95GTD5Ev7fJJXO5q7+k2KiYsXiNu5b6CdOh0v9zqt36+qjswCfEgkJxMEFvM6Le4
6FIsl8V2gGXzEhAWLBCgFABA756EUZ2W+lB4H87JaPngE+dvgw/6y3AsK3ygK0CwJ+59l7Crpkmi
1pb6+vY+4ZShug7o8FU1eLsmKzfhPpRFYTTnbRDm3kJwSzW5Of43/2PYqETqANfmwbNaXZUZDQOR
lWjgweo5VcCWsVFnWD76QMP8Ty4Mjw2q8N6CaU5sfx6FCO/JQwkp5T5LtChSTkxB0c0NcmM4ykpG
QJMSputd14ZH68c46AcotvQjOZbrBMDGYEYBm1SMa9pFxRC0UsJL8H/vqtY635n8RP5hC5ZewCNm
vmjhjD7jnsCbYdf63NhFL8gWwmPEUxIHvUIr75ER+feTHptkjCSCf5sCO6S1574chefU+DIYN9gk
v7t3jhdrntyxbyWpjduxRBMb1Q/vBBfcsS8eFlaJ0Vp3Lu1kQTiS1PEG3RsQS7c3oo12dZkmwt+h
/F0YDXrplAoXVuIG438Df7IHGHhzncWY43v4zuQepMsgSARdgEWqSeaL0P+GBrExapOt5KvZdsb3
XEQsqMen3DFWAQJJClSkauS5SvccyS9q/yUZbHzCGKScPM2I86XSMNFA0TlEMnpbEJxCylwjCMUq
taJ2X1VZO0iKHHD1xdTXU3mwwh2ZRHbO7JtZNeH9B5b+MjMR5iiPPBKXi/Y5RWd8rQcE1OQDqOWy
3ji+P8tplBXduDx2XB0zsByXNSAP7XI5eUaJRsg+AbLGH5pR/FaYwTPPF0GWOU+pRcKUjuErUt5c
K8Qj9YgD5+SOmiEBWQAzp469y48jEQL2AhIea8fU2gyCpMaR9piQRUIsJ5/I5zA5tHcq/mZ10btK
6uBGn1vK2RpbaSOd6THHY6zYfZS+VTcG8R2JVVU8BMIGgycK2ob/ZwHTmIT8N4AN3/2B7CGzQT1f
JZ+5kKetYd1gPfOtPj7357KWb/Wf/B3r3njz142VsdhxxP1G/FQKw8o6Mi1oJ9T/uhzCG/1s8w6x
SnvCSfrvJ4R2YyvmE+cpkLX50nJBNZCV686EJCA/s9DAX4xGqW436ywzz2yupIYLtN3gR7yNAgJr
09yDrvWUVcxP36++b5Wtic3LwqiT0VfsAppxgNmEBDS+UaAVHRjlhy43OEgYxSQURAbfeJQmhdPX
0RUPIRnpydBkw3501I3iyuQl9Fni0qL22iiUnYUrfPbs0fuq/aTxw+EnyBRhR6zHQKWkpJfL0Vlm
TzbzYc/taB9PJ9Dx3edyJuIMnakw4SKFtMZVILULZl1bN8d+rrgLS0pudSDf7deuvnGu6Yb3OGTf
kN2MyHDL+ILm+JwL4qgOyPi5wrZytUWlYsRcEl0jLO1Ld3XbAP8dc1+S0V7RG+naL7ARh/RRZqkC
Rdzs3Rd7Fmd4+csWEsGwFGYE0xVkTeUf8SdU3/SJNfq13cc4e6WB3x+fXYDcKbjxfPZ5YPnazlpY
7hbycBN5Sw17zGhWuxYoXHUdPbd5IbugShqCxrjFS/429p2jPhN9dYik8WqfNDlhq2pQQAaUW2g7
ggPo4slmlXBHIiLTCXiz1UP8ZmwUx8ytSoARU3Pvb4fIwEpI2b4f4uSrz7TFe1GiHvx02qzSUlmp
ocAMR6TJar0WtcfLktNHjn5xEvP4/eSoXxS+Gr3jVrxGaNNhvpnK59hwhNWpJu73mZdU/RECLT3t
7DdJGUf6rDmSxO4YTFnNzzlpQO8KJYefuw2ZUEtDbEpOK/isudbbkZ5RV/XQgZR4OUJ8toudjJPE
NdkIacDFOfwmLdD3BPV5QHueXRgHKNzrCkSclZ+ZT67jDeWkc2FCOYP22RqAmSZLHkhqiuSJ8W2f
NFfLQKbnHTcBrGtkE8r43N41gRL3QR7UUMQ93ebMgXiLdOj1I+Mihf3Q+Gx738Voi2oZT96G6qZZ
yC09jH3D02wrp4HWrYzfE6SzObZsQCaG5DRhuWcBwtVuP6Kgaa8WqBSmJ9HgW7sGgFFvciniYMNR
0KnsTLbgbbAVoNCqh+JLtU3nPWz2fDM0Qy9a5yvcmH2jKklpuKvdBrRsv3WTVgcolGEH5j8dwI7h
wJID/8mm8g/Igiy9jOuZlvaR043T01KDExPH1TT7KVaL1LR3uk857i4fS4wBwght4rjs7hPSiooE
XeFmDARjAje4t7VnqwIF9pDYhxQpOM7NdzfePrWWfEa1RMwjto9oRNxrcvF8ST+UFR7jJUQQWJLl
zhtv+moq6muev8kKlfyA8qMT2KqFjoP4FUwUM1O0Tsy0X4xQ4BJVvadtWwNEqjsJ5uw94yr4fHHC
6l3vYXPVxzFITctbll+inIHcNYNUFmK1LQxv61XiFGLHBWSdQVv6sajzK6kny6bwRBiRruSdVFaR
7DikN9pMU9C4VHSGxB3gKL/IhQ+hcbek+wqqfAPaobuTVXlYm43I7fA/eqUAWAemS2I4sU9fj1h3
Neh1swD26OsaQRvwPNiHN6YBvcYJexSDVApT5Pj28MsSK2fOOf4+jXXZYGG1L14zgxPeZRuTUjZq
0F/oLJV0iGGG9BOOhCvFBp7rt7DEIcrADM7psfh0j5qQZPZK1M6mAsUzNgojI2BRpNCZpt5ahq40
pVXt+7GMce2U/Yy1DSHzQHNbaj2CRPSkIFbc3s1QIreE51/G4cNPcXfcoaG2eo7NFrp+PBQOJGFL
+D0/N3t5FLjmyVvXOgZTFtoWalxbM3jSNgZECAJcFqbGNEUxGXaIhWBNq7q7SnnyYTwZzkn17HSx
0Cqz6+dHpV/10fz0k4eROYukJ1fYjExaJ3cjJuDyJ2yP53Iq8+X61O/PuoxejQ8tqqxw+L7IHTIm
4tO0E+lFBLanpBFGnckNK0qmNAaym7LbCrCBJtYNpctus7J2cYkNa6ECMRDaf4Az19Hqa/3m4mYK
bnVkS/SshgbBkvyMGCis4caEe8jdoEqdFHZan4wD+5ywt9RGwajQr15rdH5Zjt2kWqGZXwRtGzIl
vZ6mWQfbF3jFEknbxrvUteJvkBPSCwr/pwcMCzcJx3lfVXk69EkKFoAbPpdH0WGTv0aTJISR8voW
y5IiRWXuZgzoEIl5iC2Z7FkcyUZijH7NlQYREUvRT6iNqhtGzQIMcvxCKkfc8QC9t2Ja8QsCIDGf
xhTQmz8gLZbw7a5Q5QKDKbOHU8mnZLh95hhWLIF4r/RQ2JunVOwq1k8pb72GopNBcm6k0RvgKZ5K
AByRu1F8fGrVdhe5ZAJEizo3KlFZr4FaXA4Xsrzka3W4zxMMWNGREiGbzK5rjuDReNYNpSEC8Piv
cD8hkqbXgqckkIuNbslEq4Afmtpv/mNPPFjyiklT218fAbsTywlFE8u+g9qYVdjhXBv0aSeWDzNu
IA/qCInYkDjdPhski8Eo6TYW5OyzU5AM+p7EdN/UOBo7Zlla0IlrkabZxJkBCyu5zIfx6URx7kkm
LDymSEOz5KmNIlseLr0/xeCA4gUG5GucPfj3fe6DCO6H6uBBJz8jcAFgw4NmOPfCrrArBXt54TH+
DrOmFIs1NOVUXWBgOVoBXA2icEe39H3k3Hm3ZD2zMDhoeDyJPiGKXUgXsp9melyoI9M1EBCoHhgP
lJG/m4mdt20wcOiVDvFKP6VQN1WxuPcLoAjlTwSWcFgtRcdw45u3Ye/v7yMJFqV3Rsb3036nltNc
CnVXjYqRMjRkn1IGPmTBdl/8G2PoTC5IJanrRnjOPifeaC0b4IkMS9qE0ltlpOybTrgpV42rmkUg
Twv5+Rwp0/1rTNybUe1CA52v9k2iLDyUPOGTGuLLTgRnW2xjEm8VejcD/46CGOaCLYSGmlG0WpXr
ti6QVpYvGim8uSTKq+qrzBTyVizt9YeNAgrSaxfb5ifYBJW3a4BKmdnKF/4iOM6jicY+oLs4ph8F
2IjLCls+KosKImhFHDuHLlhQzLtKDpWwpQGyQ9sNW5TNKledB26FtRlSTj0LljJqL8zMDvabSMSk
ZChw5oikdd40G0LwzHm7WmjcoBIC/jeoWEEEcj9zbpjz9I22IR4JAQJisFCC+B5GGpOaNvSnS0Pi
7/1l4wjThcB5MxlzH0uycjOSjpup1EEuVX67BbDGhMfz7XMamdRHQeClk06msjyfzgvcPvPvAzEJ
vVvS7wnHUftyCd9OWUwTG9hYAdNwteJgGVDp3soY8QyIol+gfH4d29wWiWzWc7/R9yfN+siVEQrG
BdHOfv7kJI8JnViCheSA8L+NEoMY58B871azhy+q4NpQMv5q8sqdwOkR1EPyZyBUA45/Nl/k7xC7
UHfV5/joBwFosG26nNeNEvIkoZEzr7ZCgHS+Gfetw78TqliXYxli9IkUCoUpHSFJRQvwJF4FDmOb
jeLoPYMdhhP/rzs2W/fO5/xgIT/g3Mh8RKnRYDbUoX/umFohZ7VuNsZvcNzyrKXS8cvkn7whHwgt
+vUDstSd8sJ1YXXfQrOJxZ3PWtQF91qUOEEjRcClaWLjtrnMnqJCcQN2eByQwNhBhbwJvy+r2gbw
BxKDVP3RS41osyBdZ4ariKmsqM6cWyjhs+glLiOuJkx/5Z5qvyqbjHTXOfpMRHvtDuwfSJZEbLFa
N+Mrv8r9Wfqm5GTShkjj3adUBPlyEPky7z68eVEb8UkY5hlI5Ej3UT++bTdy60rfXY8O299daDkk
giWFQ3aX8M3s7/LTZY2z5Ona0T6XVbx2w4lwdalhyOb2kq0QfWyZexlHSbejZHRcUiLCX1v1ZMnj
toYcnzklGdFTMhPZRvLD3vd63WgiTe/poUnXNPCfmDFA48aISBMed/64lztOMz1bMRp0c0FjYGky
0ZXYrdfnBUBQUhBkyIz2XCubaDgg2Tsgj4g53X1tKQFF3/gvsDV2xxLqhCUq6/gBshwh4rAS1V5s
VEeLEdayHeDQhaS5hhOrdF489/c11f8MCj5J9T14Rnkm+vuZmgODpiPSIFqEWu64lw/2UAnljJDO
vmaKgRb2Kv2FaC7xrf9Tyc4x8icsiXSmWXgDxez8kOZZ3VN+NOyHdj8tLmqy3pHo1E3+k8Cwl5Lw
yQjS8b6unJUb8wxz52KlHJlWiOX3SUootETbhyBPrGL2rF9g5Dpoti2mFp57WA7/JOf5/ALprkRV
BpKZ46O9ch0jkr5GQMQEG4uC4ZU4qFXcHjwLGyyG3Icat4kFj9VN7eQgk3HE4KOai15YXMHWRquD
nfBhX3ptwuA844yTg9VYiULuZ+A9pRBzx/0xcEN1kUj4Ni65nuHFMDtpctJyMo0h0uX/qvLwWQTv
FAJikaOlIf4Gtzc0uGWj+XMoZV3NQ3jTktSBEVpvcn9Hf2o2cukfNWLWaRURuGzXJi2/pzALeOwz
Mgppo66NThEuXgVni4KpSMgumDlNgJHcWuUEOtcq42E6fPELUJwQjDNqRAuTT/KPVZ/YA21/aCGL
dEZ2v7XYwa227WvKfrmIKKJu6YbYmrtZoh4UIXZUDzup1T7C6I7Jl4tvUEMmGiQXJj2F6IqqgWE4
7uXAUXTJwD+T6fqo1EFx/Wi26dwWjuLyIu6knWj0Pm7BuxkUS7sLf+JGbmML3z0zHNIGwlKQGQ2j
VtSpZ7Mz85J0yFQtJ07Qi8BBieNWOgSbJIDwfG/si1nDjdnUGG7smNeGeZAJBGfyy3oAbVynI8ED
6ui9YV4G6cAtE4vO+mdvi9JafK4WPf2shdVYi8KbZQj752+H/9zB3MjQaL3OYqHwUvbXwV8KylFq
nj7THoqpOlB9uFMskuIjm6SbJTFYubhtmxGnW/nmqKHAQIbRfwQtjB+9q20C8WC3CGmEdvX43506
RxF8rSkqCJ9LDFu9yNcujjy8cuN5Qk2eblWeccegH/b66g6/FcpoNaf36InKFzVaHv5d8HY+fM+f
rkeqKvT/odHb6xEdeTZLvpMM6xI0UovELUhjEke9zDSewztXJAog4elW8dYsSAsA1JS2c8O5tUEW
0XwCUbttJyo9j9DQ738EmZj3mUZdNyAsHkR2aomeAyQLTrqUNWNCajb9E9NFboHC0SAPrvaumcQx
RSyAAw/kiobg4tkz5uIlpA/dFaiYrMJT2l2z8EJ01tGKlh4W1S8UGXcVgw7lSXMmmtdExv1TAdZw
mBnxshAn6z6BYJCm1h1bxInhHDusJ0CH7OwD/NGAavcOxALkuQ1q0Y/Nvmon/SLbDLytiARZSpRn
V1SkvQabQCQ7NC32Ibl5DpV+4O1ZaXd0L4ET6i/6Wjtx4Q33BUp50rFBefpZUHBRS0jeUrAPz4Mv
4yEfsaUhVbuNzvSkat4xNbCePlebcZ1rmnXJtMbPjvbHMOo+QKrawSsWIo6Gbw/cgV3rN9xIQiZF
FI3/v7Fret3BxDohBoCs5HeUGVAbd2Dn1z2kDF5FoqPN8Cd0DqZiLc6UAfVzEU/tYF4fBMCo+utn
cxqu8pmIwfCLqWW6lTwxGqeN9GLiRleMX5cgN/ffiUMTlL3SWFwadwDEeJCDk5AZRBoxqAilLh+J
fmqMiCsg5ogW9sI6UWmLs21F0x5XclZzvwdDUkTlAzv78uPkWS+T52XvwE5Kw+ClMHruxGqSPJSS
IZgqOtl42FZrvt9UfKoiJSSxXdeH1Z/cEDr9ww8k7tNXgFO7T3xtchh7Con2MtHC7QJq5WICh+za
7Wq9JRQoLMVUBHWIwiz1J04BvTjK8rQ9LFRnAme8F7v47h5seleRf2t8Ux9P8s4UKDRUE9XaOjnq
qhQtMsxA3oy0HFrJ2oJCDzQGjisRilKg3P4ERilx5DwjS3SZN4eewOrQNEy+3Ury3VP6WRIYROhZ
LDE0ta1BrXpgk61ImTz7IHnaRWtrcDb+lLl9U1kFuOtAoOdUqokSASQ9cszpYSNJb+GDtKKkH+gN
i8KOjtbiCMz60R65VHwlZG/y17Ejh4ZT0ssFEjAsFbAmXwyq2Q+4HRmRt9S1zS94/HFfVM8y/NU8
KcxEMdHgl2Bx9E9s9VigmD5a1UpIsLsvHzlTUupdEHwPo/+DMxafHBwD9nVlbZ8nxVrXLmqrkPfc
VLN+bp9oSZ2KmZD04Tpfks2iuvelalhjoOxRsYFwBqLcMoL8jORqXSNGyKyxDqrTMu65QmmyOd2j
u97VdOX7YN5pN8r8ontDWmMIwhxaRMB+semU3/VSRYmGd1EvLjhEbclfmCKE6fDF6sEBy8IiVeW6
tkPGUKfRtBQmUAtQACL4iNlxK0asAi5KJ8NaTMpsUK5ZhR5pvPcCxgxnXFmkM4x4Wm89QYRAUcma
IgrCXIWZ5ueBnMOXv/f1iuobTESQ2/bYw7oOFlfvhuLImukr3GgCVq+zMH0KiOKBVr3ydoz78UxT
8/UsAJizl4u+zpc2F0HTC9dABs+ilLWVkdbrzZaMxa7/g8rgkJpTtVM5qQE9/FsYiCqGA2Gb6P8r
/kDfPXNmPDRWqYMfCjfijPVmh0dKXZfVJeRhcNLQ7wHa3bnZVPSqVT+jX2G5/N09zPhIm4QNqAIy
jYj7tyPjbOwsxcot3GYTZ6QkTL/pOaZ2uXH1wWMTUv4CY1Ie25+cB6tdUiuhbYAbQiD40dqU1QmG
1HARBhh81GEA94AAn+ICjL3Sratw95K+nj6UYUop2ITuhE/XzJPVGM3V32z+Tn7tSAv22PA59ijA
TJAoISJHmaXLzhMG07DVWihlKVQ7KzpVTAec40FPJXXjvKhbENA85JTTVktIkvPcVM+zbUM7M2xx
zPnuvwn3MXw+tkTblZy8e6yVyNybFCpzHP1XTzpQVdMf2eyqcV/USojBGFmDt7hg+vbOqbx1l6aY
mBtL75OFxauWhZtW33No2cLU72KPqyFsNPFMgGuPauQe3nvutXPGPx5W8sMe7qvNfhuPrjWDoLuV
NP1tC6ImAAgJFtNwRxSDmuw2tGpXsr6aT//ivOBS29BSOfDGrIXBCYxEUodTei520npI8b6NsCYG
Gi30Af68d5dln2U1oGX94cUyrmrTsnhA/4/dcJkoE9JXzw+wmAPH8sWh35PYYtw9pCvtzV1FFrQ8
FFvhBWhMByd6igN8GYn1QIyjZRE06p1LBcsiH1wYPhuEFmgMEdX9h642j9KXE2sH+RpMN0BBz9wC
sMYGZ1K8UxybolasqaoR721F/RKNg5MrbzQxhqlRj5po8J6FQiGtKl41Wg8HdU+JPdr7bsjLVhm/
XRl7c5rn1YqkRnzhUSK5OMdE1lMhEI+2/et93zSbGYHhkzeiUADs1dFK1JY7xF4vYwQvzi1T4bMC
U0vaQs0T4ir1ezotk83xP9vjGqMmJPxrUFhmxPqJQFi8DL81edEBhKg4redh/T1OylFwvdMgXsZY
p/2a4ZRY017sge+JGpH/hH905S6QjH0aeNl7GvtQ9GwLtR6+S7CFKwa5eNM3ec5LvlQRlICpjoek
Kb4WdattiNHMloobckK4Y7Zd17FNUKPmDwcKSAn8kMvK0Y1GL5s4B3lUxugSO5WrkZWXrwyMF6Qz
OZwdBLLROwLeajebKmrINR+POd6mE0KOpPB64AT+gEokApgMgjchKEZH6Neg3bIPd1Jdq0a4wtyq
T4CA3nrSJW2Kka74jKd0ii36Q+fAGbpcPMuW/+4bSUy5YhrnPWKokseHoRA6iXCSc+EJAYB1cnqs
IUXnUuEzPkrKaduYY/C9bmlfaR357pXZ1k6H70FW+Uh+tWuIfQsjWVCZXEj6VvAqDCWPZsrwBpEJ
hH1IjbUkpv4JLiJkWxXVNOxdFC3ZwdNM5udCJOE6c8EczefRqrvN5+vthX4YrofPNQdaKzXsLMPl
Gh+UKejQfT4gV/hPes68Qld4hEKEEiZpqrnsO22fa//wzbjHwf/N9b29bN8DEMGov80VMO7omVqs
AZnECAXsDAu8jFCbIopsnSoKgYZ3VgVPD5GHe6WWw4fBJFPPZII3+BWmE4lonR797XSr8Ibp6qKF
CWxRoy39bvuFs1BUBfuZl9mgsHdITAu5I+Dx98xwXjP0/1eTqOuhROcY9DQpgVZeLLHiJO7U3f6d
D90ewJ9Eb95NOc/TcdPbDzPR/YwyuVHi2KYTNu/vHbQk7UzuOffe+WUyKMMqNN3JX94mEV36lWuv
dPYxvD5oHeSou1OunqGqeZyAxmEM/46iTtqCPJtG0WU5E3LiSnTdnSXfoSa///AO7bQvrXrc21QD
/r74EL5oq3rASCf+S0PNca/iZbv2b36QNgOopEw5D84aNwEGaQjP34L8Krg5V79YMN5/WfiSIqXi
mCkC4qxiR/sCA33bqnBvFntTX0zSYDX+ZlDx8bqLMBZeTz6OpJ6gAUwUESuEuEO3UAQwiaEbjYLu
EszmT2WrQEx8iOyqCg8/Niu5Shd7VOWypW9GEyIkhsKriv3jLfBoEMr73ofqfM6ynAwQi135aZI3
AWkC9Rv/joPerM+imBwLxr0VKyFH46CulqA/rxq3o48ziR5W65G8lLZs5g9CO6zaSnzrBzOl4PtV
jwAZpe19zY3Q1emE/Iw+/wnUgTFf5mysDxNtVtnqCvJ+3Ftdo4BFbOLxedfKTYWJy97kW2mldmgc
zMBIVym8zxvjCcoZT1LZoZaR8enZFkYAp+7jsCTA314StHcR+vMEe1WzGxwQa9xgiMnA/hUShr6/
//v0WTBB/ycEOuCaGjhVlMgqyqRhpIbfeZ1GvAsdRmJlBY/73vm+tC65AU4On3rixKaW1hnoSr37
3M9gg7Ed06CKuas31nqPZafl1c+Z+1IcBXUZKUU+FEZaiERSToM9h8UofKHLYW/cmyXXruyaGpSL
20refyE/aDU9TPwI6Kgvb9ZN6fVDBTxygAP6DawahfbICH0spdEEhaFaZEcaBTxaTFjlOFoHJ0nE
hCpVdk6DzhAgKD8T5pKeQe6xo4Nk2X3atPS0Jb+Mp3e6pJyIu879ER37YqkSznDigvfwOLcgLlaz
0u8X/CrrPNBvtvNcbMw60U1om6U461br4yqkcWgk6KBCkX5FIQin+LPvKaxysk6GTKsUA8guojyb
PywouhOziEOFldsJtPYSknmSOUKEhCHL8vo8X9BEaWlVEI6CtYxQ9NTj1CsEWnMnx4R/kAtlw997
3/C71O0fxW2cMet/7ZdijPWskXMglquERbXFx16qYrFuiFigNwvJbCFjS/neeT6U8MCeYoWEOLGD
kaOC25FiERsv7F5H5owcnu8+dn7Nwxz+R9+WdskkVwncb4f6h6JPx11t4ozxe4kWS8pKIhHBCRa0
+yXSKNvX27amXASo+UoT2hpOXElF2lUfD578nLC6yB2+LZ1XxFJP85ahccOVbpgmS5q19kkex0RJ
uIz+JL1wIqFWgpGdUWyoQFLXvlmlOAADFRYXf3gVzUYGu0aQJkjd0oAql59ibDRLq+zlAX2qKcSt
o6+RlfGOzw56Y9jOwLbncxDRBgHI2kJiBzkz0cBAEAn8gDE2cbtifs9kJ5fp3yDNdS1/oQ9djZ78
SqQnUn6MBaw8c+/XWiWDtCsylIDkrU9n74Suf9ipL5CU25EFCdUVE/izygSqO4BRrcxu9JXPyeUr
IU7HdHzBFG3O8Kj7wxvcHLFB1UFDV3l6WCBL1fcbvk0pW31m5B4I9nLnU9SjSc6ckbxQgjRJJk7h
P755dCg+ELZSicxGE/4Gwi48I41iQhtjszSmZtQFRpTk5e/89WBiOaAk//m6LYrzJn54hG+ITMvo
K7BK3VVXBmJJ6HdE+zE2WxE1THalWXYkTZNZfHhHcR7ztb5npAnpj9R3HXnjF+wM79pyEJnH1xUJ
1duGdPoxWrSVE+MLT1BKO87VqDOGt5KMbZcBNvVK33djlG55veM1VGq3CYv0QkbjPHcz5zTcbLNN
GE98zv+JQ5rgb60dEcujjUrR/OnCJ3AsNnX8siSQqGARYcH3PrbNmhR0iHfMMBRkm5AICq+TM6fB
PC2EUsA5ks1NvKFPVEAiZMkh4e5uyNbOqvwy60WcYm5wntZGoetKaFzfSFMky29T5xmjMLK9AZGw
nSXmS2T2TbIjkUKMarSLABf6gmkncZdeiMYDK84Sv72pko8Jfi0qj43HUkZbGVSim5vDIYRM6BiX
93k2ZqRqpw+p8INuL5g0mQGsqWSB9Qq+lFxXnx3orpPaZm67R5zXRpAHFB+lBRenW80MXkpqdgHd
PlZrjL51gdPtrU5jjjtNXvTXRTNCmBRi3WaWhJXRAEFnG9rf6Cnwv0407yAHO5dM7uQ33AV67WyY
SNysyk8ardXfXggrWIZRKB5jgXFVSdfIi9/IQ+W3jFBeIpnPi9B39W5k/mYEdYq56yFCeqLcPb6a
l7AndPnqxyhoVDahIOepBOv5P6dT1zgvixzgIYNirLLCRyvIBluxjWip0MLwiFMFTUzJYkOW5kqA
BTjH6li8PkHY57I/Yy0ky1kKHawdByLpO/xY4PZThnYpU5b4NorK+s95uiSRCf0z+mjCswd/7EKx
Cs3vFT+lST2Wdor+4vJu4Xuy9SeTKL7IHvCHB3jrilXVSCGzTrSTYtBYLs0bUV72RdoMtUxxHuxI
pz6ZoAR9ORgSIh8vrWnzRHMr20XbJqCK731TEmFDhzAf0hjmUY56+25HgJZIPPQ9rxqSYHHILKbo
8RoL4/EHEcRH9QovWqUeFv8rpz6cfJpMefTGoT+4UGV3K4Ml6XGMH3gv7lFtH5ThgKmfyMHdxubI
XEGhH2H1l258KBsZxAk58y/rRTUypwb0jVDlEZdVSZ4s9AmIqn6n9QqIXG96z/zs8xI42yT2ULvH
RjBgzHfTIHe4oliU1ECy37O9iZf/Wr4q6FqhPw9jJaiHX/MJ0U3u/H5i0cFAtURZ84g6WZk5W1J/
lSd3MC9cXhrvLlfFWmcONbfUAkEcSC1VQJBKapQ2Gm1b5BX4H6FXpMQmdboykJcKv2ppgHp1jKcI
DjotYBeUxmgWbBA9gXYSmxGIInxO+CkOVYf7dy3tJdW8wgRnzd/C8rG7nu/Zp3s9YrA9ngpifbQZ
V7VrAsYP+sn5xqubj+3t8NLkP7Qjfivxv5njVmBsf8NfgrgibUnscMmxn5cp8axKGtqeHpROhBry
QiEY9fILhaiafiVceV64/GQEdPwJjWqVUvBPfKIUPxDRc3R7T5yljR1l36Mjq0EJ1k4bG3WaI1Xn
1UCNG8+fw7pfrb8yzBHwFgrQSKcDMGEjl79lpw3/JHMQvCeaENqdCgqtC3mVTx1rWE+Mfzd3ke5S
6Aoz4vfZ7Q6Tg/SihWqPO3f+FxneCxQFGHVyhaVHlNaDOeLTvtrosuZ6ntCui23Glo0XfBT/tMsH
zV9tj4Dkdn1aneL+cpDXEwMEh+yuA5iWyf0pElZC0sl5rBOXZjsYnroVqGVfDf28NErc2Mw93sCx
oxhquEi8RxdawdbC2dBXIlgPULN9/ZqnfexctP7NH2GeLXwrKCyKukSra0Br8CJLKbBIDI3CYJj+
PHMqLufITFqdtaRsix5Yf6fr9tuUBJvZvy3mZx0mXIuU7Sjb2ZKfQed+Bh5ysDzta4ABhkwegXEk
ALiS09UxXMfeuGNO3mcju2VpCHkTbrHQGC7y5Xv8gXKZmpvVlB4tHmZ4ea2BuYELsqIC4KbXSuMm
rDXvxAL1E9SIRUOu3mP5tLWYMyD7ZJ7WqTnVXvFc/WslkM1kB6fp/Jx46IFP2+hPeP/BEfp8MxeD
ZllnYBzCCor3ETqHSjaNBkl4O1INPW+99vtrDxSpIZkP2oQ4H4yszYcOdyIHPJZCChHE+CP4nCkc
yS+X5hIkvPK4BhgrWmVfmQHxgraQrceBiIRpwJaICAWI0HbXHPoWhHBI8XWk7yx9atbExa96k5Pk
/fjxXxhEka1E7lvnZjSqVd6xhe6xMZGMmdMY1VEWo0ejdB3osyRdIncCkd3vWn30jEh/FdmA6pDu
WX2kwAoPVYUrmiGaymbAwYT8FyWXAaQXz+L24uyyk0gXpT6bqkH0mgrwfqRrxI5iULNVPSZxlMtX
PORfPxuN3B+e9IaSmyH5T3CbSCLiL/irqrYg1MomPUQAK2gZXWTh+N5u3BnUrjhW8rD5USKAGyTI
LcQ94jtyKnVv6doBgb1v27TCgy3aBE101ejc1ENJDRMzBIhevqmAx6lb7N0UeDJfec/+lnOCDfS6
qAp0rO+EIEMKg07dURu1HcxsHf/9VrAqTDV81aWJD8++zT78zPb2RQWxHRP+K1etNI1eaI+mG6U5
cfiEs0TgPvsyC+X93jPlYzHObPHl3kAn0kkFGN1DZxz7+jbvUAb4bLYNBjXDxVHNW2Vwrp86RSGA
KaQXPWpJL8cXM7xJipFRmI7/hMsSv4YJ0ATbNfHo87fyE2o5k6y7Cq0GIduQJW9eQat5CWFFsfg5
7xIMj80hJk2kDpaCkcmje4n35Fh8bncSur4jOGDYTI5G1Y5QM6arRk0osmZHj5osXy3USGs9AWQp
ihONRNYSIEojisrG+jrYzkEN6wJhyucdQFao+szoREBt0UjLzbQS57IrLQikzjURqVv1bNkK/ev3
nVhBMK6WbO+G9Keaeqk3epbSSmw7cATc0jUQRzkOkIXLE/31bxPlNhtMnMhgBFIMCOlzyhTjGmNb
tvjx4jFUy33uT41e6NBOJZ9P3IJBbJep2L+imAy6YW8j0CEsub5JXl8Ywa8Qy+m3eVULMBIZQcYo
DUFsoF1YmTC9LBfIFptcvKYsgGewV+iyQi5Fx2bxEY/Z2G5ITQcoNWj3ODj0nIlPmX6CnbxU4TwE
jolqSohQN2LWbEIBtULh2c6FY+adwUMDzAKDjMxxJsrbucp39Wyab/9Sd1V/3qTK3bvJTZxdGbwq
KVT4AHDKMdkogPE7ma1WBc5czRUeW1pqHNOWaz2rQG7H9Gcex+Alq8U+vBoBzgy/ggifZr9a9hrA
pYZ2TSSKkTAdGOH6bwPUKuCK0BNM2mtmQVUFmojXVgV775IvDHoMrMCGfLZjcJhgwveQSQAbbNzA
83NQpRaXUo5caDEPNvQVoEavKhs34LE32fNAv2dx3gR3Wfy+4NBy349GvcuuNsctXBtiVzJGK833
ljKdNgYkt1gf59hmu8aTHDxt4281T1FKnMz4b3WdWzszk2fFmrbfK5NvX++bdKEkk5Z6Ewfsisr9
QMEBPt5meQxcGrX+RRB7Doeiz0LMgD64DC39FErlY+WftEBP73gk25ZTSXiKNMaO9x9nT51PWr2R
aeQH1kWyIdkpybo/SnH7bnU7Iq4c6qWqhqawFrqZWLfrvCSVxngUFwTc+w5w1YIVn2AGzXYDun7n
BgU4jYmZiLfAtcbGv5Py4dW0ogm3ZHK217tLrDaR6JjU+2bYnAI4vvrlfoDpqcld8iPXU9R/Zb+o
5RbgEsb/O4XwIiB7KjqWIbLXA3oJOMhWuQllUGfAq82e9OpsQEhhlqoYHHRAWJwZnQUJlvc9Bz7N
feJhFqW2ZrukvpEKRCPYtkrztH3WCvYbw5eAwp4CFpyCiaTzVuWWh9Bt9mhAp5iDVVbZ0XVE6qC2
nzjOcW1NeCgffbr9dLiA6jZB0Q0L3um7lnjLptsqB69GdbxLEanpKC3Qhhr5KxUiZr8VJFGHqdha
QPEKDkX0We+XSnbw/Fz68CN2rNC3z2pgwSlYXhHtUVrv4aOwiHe56dECtCilKgAb78g20fwKbC4l
XBu8aRIQ4WJGrhTCke7YcpEi+n6EMsvi90QMUg4slHyKLmavPXbC2PhcygS1YnQJTwPtmj03/3rT
ImSo9P+79qX+rtIVq5ZuImxuQWL6G5tY5K3edSWzi/R1GeZO4TdlbqPhshMl3K9FlwyWo+f9wsV3
UBvwgXLL+byvO8XAMXvyFrbvSaQE3X3LDIeJmpmlZtbpemilh90xu95qdGkAZmSFFrxFyQIS9bI2
N6jDu3Knj1/N2bDvM5bESewjjz2dE9SmWp+Alxj52G5c5IELiq1fCjurAvzDkKPsjYEvXUoE+lCh
gRbqgH/e0O3l+gaWJ+mIl56TrgGvpARvkAN+ZTdDimegf0Fo9z3Gn2lB/+7Ofk98UUVbGCKe77bq
oXK8Sn5pTvr+TbgjHawao5O0sQWrzIMn8e8WmdoJTalfLynGYS+3BJofXk7FPrrABnUYWXbF0gbB
XtPdpCB0p46sLO6pjKeO1Ewmk8x10I4gCnSfZntGLrvXM6FEYsPNBptMeIR7IAYS37iH0gDVqWb1
8Wg+XscbHRcA5C7Kxs/mPPNCnB8jjqalSudELH3Cl4AsAAcIqQYKAXNKkNu8PqwdYRCYUjVyo4kQ
zVvkvMZtfsbBvIhLKbDicVAU+WcL+AFjgidVckL3s8CKq11MwWFz1QP2Q+ljBl4n0xTCiGkn+52P
m4o9b77PCRuZ8GrJhUeSJwpN2LgpqpPvQScYlEnqQnnR4w8/DXg+nDPwQudDeYiQ5mIbFmHMBj6b
7pFcaNDKD5Pj7NYd+L9POqjmQVbxhQqS2wHXgxWhYZTARcWUu5kjocbgd1YyQl5p1Na78OUr3JPx
qyOSD4cZCBjpYXFsAi0DiapKs916Yn2oTXI0CL7uQeRYzfSevukvDAwwXmZDy/6VI4Be+JL59UzL
kO1vZoxugLmdRCuFWn50iUREvKkqkC0DIa/A+gXHkV6VvlEexrJDWvP1WYQdAy/FVz9AxVxP0gXq
2SlNEDW0cpJCbL44WeWbeUnladF+R+tsG7oxV1ZlL+epNawMQ1THbDjzpx/AsPfOmxDEGx8mmdh0
zQfqheJPY/KFgry6c/p80X4ZyIJm32dv8a0Dyg+dFeKHEXS4yupkR4xov6pGcdLi1poAsQqzKwOG
gfNmojznprgaiRdL6uWy4BItBStsy59zcYU/b026D0Qz7ebZwj50tVjkV1AqXzZuKXiRdMAcj7R4
emTTAhLez6dsPmaGyp3z5JJNYHb2WuelCaVU4BeI6LUqnGQHJChEtLaClX8po54J67GoOmL5FQPf
67e0QB/f82pzbOVqeaAFpsxOWVQVQhPONNZscfmcaekck6ZavHkGaTXCyrJ4OQS58TmmU43vi+EO
huDNqwuJyXgEiz1482z5qTWV6TDc91bkqPMlcr9cY7rlietyy8f57pUwm1stu6pFvZYUprxcTgiZ
ecblji29qLojyXM8lJvcOBCEmzDraUUwKrzJsbqyUOcd+r3i4sFB3hS1UWUcjKi7Jx3WGNjeTQ8T
YkqtHORFjVMSCcTVRIHfmdYp+8ol9jotlYcGgKRnpcnhkOCTHmFex8c/VKPYfXyESaS9edvJytul
tq9skG8Sm1Z6LvXy4cWfoiP3Ec4DJqGnhn7sTBrqR+Y0yK7Iz7WkbcvCJoSpnDIgpHvmxJXUDTUB
roXTWPt2tzujrQjgBSsPyJ0yEYzE0dFC1YzeO10BVMsXJ7ZLeF4kt2hVV95V0AtpvXGTtW6xIF7R
jqow0VY2owcaP7/Fz4Ieai9rSyeCYHJb/BwBVww5iKlLGjucpBkjhe+H+c/ImSfYw2ud2WDjbVO3
L65fKrjIioLUchsCsEqWFidCbeLc809wVtyCNRJgTFZ4d3Or/uR92KMJiyY91tWQUqtf1n0WA7vu
huRPe5GbZZuL6/5+KSzagB632ZyokGDulcJEz5xlM7/52MTMv7D5xoZUSLllA//KwN/PzqYGoEkL
0g+SLwY1FNQuVUM1w2VVbvLDY8JjKWm0y9ao8KT9phMqSN4SXQU86qHg7w23cAqq+Kpg3gvtb9CQ
JbUXZ/IFXdXOTl7IK/L7tnxBRCviRlEdybWvdQzkhNxJ+jH4Ebw1vRSeivZ0GikR+zkuakFfPnZo
NbLUvXsU7dTw+BbqlTb/Ewj+NPS2HdC1dbLESa7kz0iwuEHsg+h+U7czZyIQgjfd3dfcJoerdYAI
MYLE+s1bnUeXw+Z8gduypGQp3h/qKOfqP9VEdtajtYiP47fgMuUIBdmJ7LYxtbHAOZRa75YE/irD
cNBrBgwm6G2z7/JSlO4vFsbE7TqdI2RMEbdROJ2qXi7OHTx3lamOLbE8BOdaKSMKNYhu8ScUmj5X
plljAsB5kiE9wvElJr+Gu/EfYJFvfDiHW1dLzg9xMZyJoZ7T9zlAi0XMSncGEjWY019QucxgYo9i
vmXEV8XHcgOR3Ta9/VCh/igLNU0eP3mQsHqiNR+QIngK7irzc4WR6tuG5bOiXXyeoNd8t22yqTwQ
kgZ7YuYTIkbbaN5lUE1bVvcgorgJ5Mua1OlJKcdRZtw0X9N/ETaVubxHN6xWJLpVd2fb2ee8sIrJ
5r98fhL3PC36JpHRz/r8lQ0LYlgdy8JPnYpYCGxq7gGQQhoR7WsJ64yrRAqK1LCYA/Jo4/+3nav9
UZ1AGrhPUGsYQnJhuJVGaiwL8U0dezhUTyB7/xbC9GTdJU0TfAlKPH+voYYM3/GKq+cxw455uuvW
joa4TcvHwHCakq4mD1BgJujVqOVvrTefdRNLh+tvTCz7aL3uUjzFQJiMQVsB+GCHh64Fa9fHyQN5
+DGsoDVedTbwT2jUUAl1KXhdWOZvgFlod7+5Vgoo4bjATWl43PAHm082yVvc1wP1d1UbQp8vNUn8
lvB5gio4gw6mpjgbea2zC7iId+W7UTIfvk+v4ePrcdpe05SJs8yzDnYfC0QxwUDfFhttuxqPBHDx
/OlFvFtC1V0vsayKNDvfMPXbEvXBI6+sxO48i6BHYEpBA9vwX1bYpE8DnYIoFcV9FkXRrLe+dkJ3
kfUSbf2yywK6T05ATL7mLWjZWT/2lc/9gsVYAvEa0/KUzXas3vgTuQOSVrRHE4diJSc+n1nlorgg
aeT2sxH4HF5MnBvMSZRmQWEFizPib2Jb1QuYjWvuX7H16wr/iarkQUJ99XujcGY06rZ14ygls2kr
cnxt9pDDckAtglLlGb2smUz+Q11LgxlXvwLxpdnTq3J8iuXKuWc8amIwK0OtjPrEUZGZQtOF8fOq
CIl/R1VigY2axt7bjRZ+bqLyLS5urhMKc1qvP/TM/xkxo5ParwFyPar9IVh5sOYQzx/qoX/UgrzV
C/OO6TcXAR5O2hBo1xlMT6xTLYrQdpiwDK3MRJqrAi6TBvmrz4BcZXDORd+abtQppem+Zqj6aOKL
7ZPjeGpVvCANRvbe+Suz2o1f7UE0/dGDmgIiWkN70Bh+rTgaKX2Kzn4cEM4igg1EuHfdVXjQlSkY
a7hr8TJaYVLCRNP/np2X+BZc0JHUeqboPuNAA9fDGlIbwNzHesfFOo69mCNur42mTlJ2VVEAzJEu
Ztmao36sOK0sKyyFfoLwi2QW/4WoGjsJYP3/T1mXTnan0WWMv2kzEglCeNkKT9si9s/h/NMqEaxi
rICG4pCZgxI8c8OdfxS9T8lO+yH83DXXcCzAthciZKFMpCd6DQ4MIEuTxt4HD5eONvrQAB2asMHw
dNZeaIRE9xD269mUbC5S8dAKHqhULUw6X5uvtg+e0m5GAIZJbUn/X+5C9y8gIRf6X4zlijvJGhko
s1D2YHbLqSFkKdggvUP3YiQ5WmgFk9tfhO7Po+8P0zs+Qy9cvAFwCAy1azSw8qTHOKQbAGm+S+O5
y0D+mJhNikdWTWDGbDu9DObcGV7Jdn7xqBkAyI8aYQ+0VlyWC7QBQzQu7xGdTpdY/ceEBkSnIG+u
Bpr8Gv34ntaOx0oAI8Z8esFj08/3E3jAvFVhneRLkJfDBEZr4E0z6pEI+rpFzxanAy9TlNsi+e0C
v/tVSwAKtt2sf4eI0w4SOuFNtUjPeC1wNwf8O+Wd3sZWJ9Bk8lq6sZFtG+mHZieEB3NLUbXV/zvd
FGGk1DbTYlu2g0lVTuLMjUGz+5oTM2JFekBeGjvI0jzPqbhBa0VCrwrp3A+pgL8rHIMd8kgpWbCe
5RNDvtfWuF/HjBL7kQ0dAYOduWmDHq2TmxrHO7NrB6JBnX16eTRJfj3tPy1LSDTjKc3hJtG1Ui+a
RZrAnY0gcbjVuQDsQq3foyb9oTvi55rpzpMFO/aX/pB3bSiVMqBgy35aPaZlwIKDhFINM5XS/Qn7
CUswHELVTIIYtzxEyl8AbxGXdt3Z43VmMVAz7LmKllUrURBshOM55do99BZe+i2jzrK9i/HQ92m3
6FRRd5HQKg+Nz/4DkdKR3ES29N526ZTpJaoVJinFqwIsQattLc5+NyGoMFGamPtBFJbyhbVZsfjr
1YsApi7OAwKTSK6BAZ6qty9FHiAEI+sFE2wMYUmTa2lBc6V0AVkrml3+Cj1EAbFCoyhf3Kjy/aRR
6++zFpjPAPsfSQ0SYFrKgt95nT2HlPggV/rcIQEX1wYyDoL5DfdgYA0f4fhoXRFU/XumvlViLRoB
/ckNeVvcU1Fa/ApvnpDlfgPQy+LZe5xCg8EGgKgbrINYmMCmySK1qqq/ruW+onal/3fw3JHgPWji
5ETT99WxTnxrjzkrEwGdfhuAKpRN2qsaL+jL4dL3RWYQ2uGTLUeJ4w8yGMLthSQKnLOXGWqdabVD
MAX8Pvwj3IDGW9sU02ZWQyaWeqtdkREzv+1tKMUj70DfG86m5rN6UkUvDuixSMey++O7dirwcCjZ
4W7tS+cVWRkOhh87f9rGVlIzMdHVnoFCF562HD3zEdALcnxTzBZiiIJFXPdzu+zJWzBvrmWXsxqq
ElYAnOqDMf5lNhVZF+4bYdqcIppdMli+smwHeDBukBDFx0BESXtUtREgj/oSzUvvFvL0QqfBYCuK
QXef3HlM4mvhOVPrq+Dac93B+fd0b1YX2ctNPoaM5lf8el9YCflqVF9hZNmhtASXPi9z/VbSE8K1
hDlkBmmNb1uI8ZRHu8KG7hKjtK7BR5wx4mhIpOl6ZUDtotlV8fb3uZHNkp9xSHljuWMu8eP4DEsX
rSiVUf8xMj8bqWvi1VIwD7XA1s06JbtU+IHTpiCxkw5BbHEiRFtpJabvt7GFKh5udpUFTayvejP6
BgurXqyMdHZmjOZQmWtJ7YmLiS8wH5pb33PdI/fG+Su5v0SKljOENm/qAuTaI3dpL8aKLUXirXWp
u9t7wLt+tYjAGibVSZr+4/4yF/1vPFqpGBD/5SlDSrovKhMsYMMQdLZAvjR7pl6PTlj7CnPYd8Lf
OwdlueplGgmmUI2Dd3OwqFwOwyltAJ1aLUFKMzREgsxHs0K2TG/7oDyNFflclpyqqLICHdjcuQxy
/2sIgtAtpSydzh8QY1mBgYD58/phdSpevDCABZ3XlDe2yFJELSY9/BwIxq5v9943e7iCRHOgVsQR
ZGrkzXLnOzWz3VusbyjQudE5koX5JnhKXMZSaGtWWxIZI66Hmc6gvV/Kg4+d9g39FUkW0W3x+GAX
aET3ofgglSbUryOkq6KPrFxPTML0OmDspQvPD3BpV/uXm1ZYQ1DzeO0fA6uUZSB3cGDQcNbZ/fT8
OZp6vAPeQ02mVoiRbZAtvm8aRJL2eBKGbQlSTVUYKU9z2sD2z+aQQQax4XvRHnaRiZp2RlQ74sWN
ENFMLIv7Up6kvVYHKSOSZeVKsdzHKUl8XOEERYICIqBeicQmvu9ZlM+qnjMG8UcYokTsaOxntQa5
ol5Jv2zaMrklVnzoYhjSkvHqHEgEwx1wi1NM/KZKDRobJ1cA6l2EpuYcnihykcxiGeKT34Sr7Kxh
G6qWnfnkLnrTB3MtxCw5lIMhosngER4QaOzx/TU9tS3cCjBIEWWHStuw+RnpuVmVLtPmehg5J496
lkvwm0m8Wf5FAqp3zljnBYMGy5Z0MEKQjXj1Pkd+aL63SbYb1tVEaAzHEKaJnDQQ0v1jXtScp/jc
VdVcImBqZMI9RK03Xk346knBiT1C+iHEpLVuXCLkoQ63xf5/toPryXF3HvmdYuSQ8WHhKUKe3Px2
Ss0JS6kKpR5sVJG/5g//6Dt8tyNcHi/eaV6FpvXtA6UgrsvgyoObPEHeZVcIIr16JW9L/lozpEEt
xokb6iEugHE9d6wf+D9fwvormbCF5LbY+R9/zyX0ZcGRLk8dPQRYN8xhLi7SPv6Ggzf83h5/Q0uY
uL+WKOpaTuCxFJAXOmUfzj/Pbxdq5ltMZM74xIny+XHVHSXEUrJTEZvh+fsMrKg6+rAfdTUva072
CbNuuLf1A5QLEHBQnjOSWNmm5mUZJaqWM073MSURlo+9hk6bDT1Cg7pAvhF72X8Ce4UhZTePwKso
a+VR15+Y2MVgx4sDDihHIEZ1OERyseqWtx9wwgFfvhYmzuvXTcL5prZOIvWeLGUf5pQRWBGfYhyg
fu9nM4a2W7ePWGr1brZXOhUgtZbk6d1TCXah9InXm0/u3UeS0DxTckjT77FiH5woacropIDb/cRa
e3YTziF6N/0p8sQrOF1dPnvwat1Zp9ourIPag97YQuKiGi1ZtmNpuEqws8gMkp2/iK3uhc9PaJpU
bf8uqkqgN4tPt01B9w+Re21sxNa5vNVhQ8NI/pgVrgeL7y0RQ8SEs1oKw48h+NQsUiUFyEMH72MB
tc0J6+wC+RRgPwIPZly2qsyswEJg13uf8ACDeygjvnywM6LG4O58kvaOD/o16uziK9gg3EtHWCKH
IBDJbxhCIkfiQMA1aqogXxu8ZqZDSEqZPxIxw1uiAPI1C7SWSxInv+eHkDCaQ++G5W4uSUDhSMV1
F1b1RD+vqmCdvJmHVSuzEVwEAdDKE6hmoKZNZp/0V8l/puI9tW6OhzF+k6+0bOGZvNNiu+XqYEib
7qQ3GS22syJOiRoUwm5/80LhLcfHQn6s2IM5HynPp1YtiX5tK4QPw2MkPHkjIB/ghQH92p9Lqz6P
oyYzORS1MUDp1uMnQngiVNfQ25uWa23siowAm0lEa6eObMUASz4JfygviSL/Tr7wRCgZZjwTlC54
vd12ofJj5Wmb/bJsiCYNUhB82zsXY5HP/I2co2zJYpXxwn8XKDJD3pOLT3sLLFIHs6fxsqqECRUz
3oRS0mXBOAuoi7bVY3aWcPjD23KbgmLPKlQB4DAfjG3ekTz84CzHCwM+DwzCnQ47wlBFEB5lNM/T
FLgp0wR6Q/poztiY4BNAa3DUCpRu7p4xGwmDoVqK6C2rJ3iG2XzRlUrXiJn4gsK2UENlNR5QFR4T
YlLsGr/OUvcjlleVrJp83+9A858W5BIQ64ub1D2c8ZDIjLC/AvVpsSEb388BUMpyYuh6xKI9YWsO
tvlghPX1RNSjw2HIYdKqo1/jfOMzVS+U1IUHO5oCwyCR8QpVrWm7EcSyv3IDks18ka/Ot9lr5Qih
MVyTD8CRqdxgDT9ezd9QnWFOGa2edwqn5JNKBwQfekRI+kzapWQsIbGJi6cDZ+8iPHunOuYJlEQy
BEnCudjjXbFMgxPa88kAjHUhyGgOOJT+klkE93ZZUs6/7pxw9Mfu42p0FhpHptKcL4c+iASCq8s3
K1yRbLoEK7AwMI+q/NuKhygUYkTuGuM8yBaEJfgTKWYb5Ti2t7DxVgfKW0K+FWhlXOLloBJL1lE6
7t5dnlciXyXJPW6z4hgakvGR/rTqdmZwZ/8ST1etxcOMsitqVRlUwv1ihGMIu0kmdm52h4TL036X
NvZqN0RDkPIluo9RFqCS5Fd34tNzGEUmAmDLVG6WBjGy+uHjqK6R4MQxSKVh//i9iY1bjZHjJovk
6p8vndeczQaENHaP4gJjEq8csJERadHF2y4Z9+BbcX23ies7Biao5nWEC2rrM0Zn7wgNEJF4w6bE
Gi5hmTRuch5/AJ4aMDMc7kCCuehSzra5xsDn1RWdMZk/WZX35DNWP/X4nu4hoG5p1mJSlvkRBKB6
MnXjYLswV+YDqow6iDnM/QzttEKMFrtnnTlLNX3h88uDcNbb2Qd+wbL9gclHmpv2fuqQZJJDvTTl
+rNGCfH1nXCdhWDk7NGIFUoODNeKsxewCktas10PNcmoHnTxDB2T42GO59bFoHaspGDw/ZyNSByW
PIJgx4EvOTN8goR4o0y5QwQy1xyYbws6SbnyjM0unTuKYnVgb59DX482Sdu2cLgQHubv3x0Qgmz9
wyaoIjjDVUEYWw9Vw6qhk0BK1hLBb41T+jy5+wgWZlFD5aMvDj5IwGlXXyNg4JeO/2scIoQ6L7vk
1/h1+UwmcCzO3olO4lZt7ZaAKR8s/9SZWMauWOsbvpg7/1o3o7YnwySmVEacb8u9/sJhmuDK/qpp
Q9IKkd9B1iRv2reU5dXGo/WlZAZRTxwvXKUFqnu4LjBc03nGbSidicslChZdA/bI1kiJMjLd9baE
0BNnkOIFA7jye/qKmCub4UN6QWlLp6b7FWmxymK55/44Vp1z1v/9o/E9r8gENg3YucVgxRLCVX8f
NkNaWB1TvbZqSTpMO4cRMttRBwreA6I4quLSZ959V338/IovSLKMbUyx/moVU3fnISfJ6ZcD5fIT
fYWETcAT2VEEvpad2Ee8D4QX8Cg3xz4NQQhv9efPkyMeh8vrevHVKr7kOvVVnhnDERGYuY/6QlNT
kCIz9BtnIatCAbpkTVxe9z4hb6NZxKL5/k4ML6Rdkyo3ztzonJGW/pu70kCUNKS5jws8RyCy7zMv
Lvl+uyoCs5vAUhzrMEVU0HUwIxmdDgkj3Xz6ENXwhfL/lUOs39WxeAf7lbARQwWeNxMkxpggoCre
a17IhOSeoHRT6vQBDRMQatMIV+KtGdeeCz5GfLnFacVLMZcNDXR6CwIMYaf/hj37lqudS/Yecf4V
ReeuBkanrBicUXg1t2CgXUUgrj6Zbr4EyxXRIfQOTK507Ku7d7bj0SKUeZaytrP9qw+l9KSLfav8
G50BUPT48pXxpVf3Mm2fP/ndgeTJaz4lL64C0d2+oBX4ce6iYI6U5tgAESOOFXF3J23j0C1X5jDU
IknmsvnYoAKvQNYlwzwIPqlZvmttsZR9ISbCyQ0HNCJrOQxCqNVY+iCBcy/zZD2NEmgBIji3vpGK
XK1S9ED3eG3Mhk7AE86Dat4GeN8a6Kg3Vjzqpj4R0zK7WYXssiBAhgTkkCJh08sovMEZvi8Qca6c
yLRxzEViZScybcUVYKgTQLTvO5uELD7Mt0wgD6q5WRkmVqRxmF84SzSdL32JdFVpUeCu77sQk8Sp
j+juDznV77ogbStS23O7vE4vcxOgTM6ldoQrZPIsplWH/9xCxut/oMLF3wcAsMv3YKWU5TyiAgAj
BUHl62GvsU6HOZI3YY7gvYqSHjnIkztg0jIQKkVD338261H8yWUge0312deQT1W89HLqA761YlwL
0Vb3wNBTNVY6eowsx7tL2rl8LY0Ngcj4jq+He6mD1HJ92df0JTlvaLAJP0e6LLTLQNjO4aiSmQ9R
dsWy2v3x2xmx7PyW0oFt3l0Fpm96Co4mFbnKB/gVGIrU3v8b1oLJLM7qW4JcOlsuNaBNm/vJELb3
9BhOYLSdRakAK5thOJxH5lRAHgDj5aX7jucGJRaQZrq72d92pIgS4kO/06GrQnBQWxuJ2SOlh5By
7NZu4iJp6YYCcJ7sq60IyhPIE+ogKfxoD4hwOcMQg1JzzHr42G1NTGZtdccttqerjFOp0uLwvn6p
joH4upttQkdOy5oZowROQLrJrdoV7HXC5yA2gJ3zByzA+3UzHQ0O86SOayoi22/hzvd9F81/2Hjm
XVZ6rz0sQVR2NJCYsyf4U8R5e4QDMyxqYs8epijgcgBh3pL27VHmfan/FCA5b8srk4Lq5KDz7azX
Tc5mFDxCY0prx8LYYvUM6XEsdQypjTlbNU7t/teTQjyV/3Fp8eZVvKA6ptv574qCrGNjbeiFyZtR
HzXrIoomxadmlLxH2hC1OxMM4R96X2Wan/9vVtuiZNCrzIhXOXsFEngBGmY8opHyKn/kFaQou9fW
t526ddTkyoTgqxqIb1FBExUVb4rQTiyy717FPCzqgvV84Nj5GUZKCyHyhJFYszjBjGzB/P+HVR93
e8ona/sIjRmgtMUGfzYbYEekuZmtPOWYGgpWoFpEq0/EW7Xd9T9xK7uqD8JapYFFhm5sfYwib3K8
vDlTL6T2K6SnhnShmPgR+dilOUXOPQQcf/afcUfE54SDgeeGQ3LS1A6vl/Wowhd6RlrJlHSvOhal
qP9XX3GIko87awrFYsOXj8YwVkkft9xthGrlcQtLW84ZqipB2v3QHCDoEZpc4Q26Jcr04WKc7Am9
SIKLDyhr4HP7Z1fhC3Lb989tbgwx1badjkt6XUVhOJqlC/NcTPT8cnyFoVDWvfIoICVpBvWYLaDW
8vprJNgtx/0S5qm85/mTuaQIxNSzgp7JvgREsn8kk02mwwtVLSqfHqgOvak0ixy4Kmh7OWY+0CNJ
GKYSz5vDKQmvOxbreTGkrMQaWTL+LDF7bCo1+MF+tkwjgJDn68Cde4t2iBzvp3xd13AXhy9Zd8S2
b0qPWULgbqXl2uPZMV/4qrPC36Iqe6793qL/+bgEOqpOY5VDMY+rozbiP9eZlmiSRmNWoK6RpHob
DdziGgfKRYc7jGEgLZOknnWGg1afljOy6IJY/FFxPUl5QqnnXyKZ6hzxnHUHOYZPCLk7FEomWN7R
q05YzP+soQJ58QW866fFyjnAqRDhxZsAtUqFS4eaSVQTKQe+whKlGKVeb18RI7mCGpOFljI4+mpW
+O4iLh8qeFFHN5UWd45BGsqTDACk5w3HO6UCj1jU70cyWZm06pgFOqkZhbzsdfCsFoRk6fDx9W3n
3NXTDeAW3QJhL/l2ETGZRi//0aPqU/pDL6nQEUDDXX3LtIl/m/D4Z6rjV3Pw/kulQH9U38e8XiIr
arkZpesxlgVQNrA9In/dTtzQjRW8O54I+/NmH4kYRX1eii1KTArb4Hz9nR+kALmqM8UzXH76rSOO
2vRvhvbjpgSlBjdmiGEXVHB0sjAYLCXAcOlmrvGiGaR79EfCwIxYFwOFQxVYya7m4K8C9Vv6bTTm
LV/aV50zu+5EBl9pFByMIqiJrN9dC037enOurU+b26lLUntc5O9hAwNhvdCM+bhmoTvPWFlAms0f
6FiivL3qL7FPfgyTA21zwtGfSASJK0pyvPo+um2pyUWuRFDDN8bi+DlbiBBwB8EDXyy+kARrnXUT
FxEV280xrrz+D7aUChfQKgLSPZWfy5G4A1Rgtk1L70Wsr2KloaxAdb7NEbr8xygzFhBO7clv04Ar
hQnf11ttr8D7L52S2YL2twc5gxbFJodvHQhJaMziisizuy/iyWHIrsIQmP5OZt6kYjr+iRuWPCeh
j5Qr9PijbcbkU1qJ4rVmpH2vSZh51xjKx3MWSz4vJJGvZhQndiMkRIHRu3Glsjo3JlOHJAJgnb+9
f9EPbggU0RNubclVdgIJ8VDBDmtnnY46YIfzPsY2b4xkTaBKhxe4NNAMkQdEcCLQaLTZYy48FZ4Z
ajLmB8DVIp9vvD1rd8butvsyaJwI1Gx/CNKgZAmFaMh31lVQZm7xxRQCgATliaB+pNkNgJgyIiLa
F9Cto46O0+vXEQaKDN4XMZaNWOliZ6mOdp8YsDxB+h9gGXWFBIlicbZFzSn1u+7/0gjHHb0ZJ2vp
luYLlkN5+yTo69rNbPG8fC2tpCHoiIiSZ3Wlqs9WnKBlWP9lyerRT0PBQEAIccaNPksCypDv1eCR
8rLxDcDBWoQU8ZR+hmXp9AacNBYEuXcdKsnl7k/cUmGBiKTW/lD4Pwfxh7IKtDzrQOICm2G/8f9M
clYxuOXE/uEpvzNAzAlsn86RM93P+Elj2HnaVyYWUSm8uEuo64iEwovc6IWCotKHCkhBWGaGQJQp
aY+pk8ZKI2SRh+OjvDnzdBjV2Z9E80DB70IntmJBvdVUhQPmtSlgAuOPQ4IZWqv7k/2504Qt2rzl
bb+uvAbm+0+EuZwklGSkgKsCBUgi4d+lCE6mChn6JwWffRs97elYDhgA/yxvgHxUXiPOeAzH3Y2g
XkxjOdsmr8yXuxhNrdWrk9bP0ENqToFDpPaj25BKw7+heVzJlIkcga2C1UEewh0WBpfWoNBqHiRt
uJEgl7MyGPLKYWnwh5kq+o6Cy0bE2eBSwqeP+OxjWmBov3T4/3M7Oi2VDNlK4Axm2RbzOIcS0lnh
FDCcGX1Aqz9LpzDizwSNTQJUeyq4cs857sZj29d56GaG0NcbXRHvk92nDHWH6vueDzuGZZrhQxjN
jpfoUpxOGuItU72I8KWCPateZ9U+lAD+sLuSrgGgofNTsPM/NTXaGz3+vDL+ESzazd42FrgLq/ZX
7JXxsddb65HGwn811P0rlfH6X6SjD49t2pk5D4EQnoabN44cSrFytEFLmuKVvuBaS4Stt3LxFUCt
Pf5Qp9X2aYOomqgRahDw6HsihjpvouTCe3wd56YOLSt3XW7hWmrGusKqelKu4ObcAaRC3ik0UfsE
fAY15q7CH38WSTD2t+8/deKqZub3mwR8ikJC8Ga1fhSyeJXvNOoY9L+L9ngGhnA61oQKpaFciQNL
AszbjJgGYJLUSZONzAEbg1SHyDCVQtckG3Kjr8NTNyoenIXlksq/1oRvWOHqZ02dxvbapQHQnZts
JhEbZ2XxvRjj2agFF3i2AG5XnLImSOfE8MG3WekRBf+CwCuucL6xZ7e9z9rDdcoBs0uNpOq1Mwsu
yGC+ErOV0l6x//tUDKAshNwXYHG10TOXaE3UK3i+ZfVx5YFbQUFvw/10mtujCBBofo6Q0rdBfstn
ME0haczrgswxXZ0CFyE0HXYoiq/6aK/ZBBiKKsWF+hbeK53Iop98uc6PWkY9lWvmSy85s3c0zxxK
l+sTZJD6Pdo76y0DGQN5W25cNjP5ZQXrju98ZhIj6iJNAmKox2zEl86b3kVyM/FeSdpS1hyrA8HS
fDuoXC272xahGFV1xAlYsFBN5OO30i7hHaLf4Hdf9eOI8pw4neRsHAArnig/9QWM+GbZd0UPVQdg
xRMsB985rabkB9xeuDQoCHy/lOtHDSjZiP79pe3EXGR++pzHW9fxve9w4oiN7/Hq5OdFRNpLwS3g
g2ea4NSKJkiI6adhJ0Pm6veWO71AmhWNJvRTdcT8dMAvaW6h5+qGlTEJs9SB2UUHyRHZhjJjIy3Y
JQDf3AOJF5gR9VZQ8MVR3jXWr9R7SGL5gF6F1swfizhZ3aKnLqCi3ZFidvsYdHxEUKL+xHTH8vQw
CuAaCxDNYLrk3OO97E28m6eBX0hQrzp++5fnGYtrV3I6n/Lol/uEG2mpsxgNsabBwRwe7ZDs4CZ6
wwj4BInLC+XyAk5WDrB/E/ZzDCEemE1pKYeuY3bPBI5mAXhallOS7IqBpmKGyLeCDfJ8MAvni3yq
LaaMHnApyLDrXphCJjji4KNlCEc6bKnOLEycw78UuFLgKS8Lup/02CCQN4qbQdDNotTJiZ/i2Ct1
jIsztYqldhXp0BmauOKhoJWbv0fRvIu/kUzETQ54RPUnamqaqZRQI9+oCo/Ks40bFgR/R0FzoEuy
JfrClMLj4nw5BD0x/JzfM12G1C467skmtV+ZR6JChRHY4EKx7rK7oIZkFbyZ9eFqHFAbvflO2iwL
rGOOnTGd9z1Kd5yFCrMslH/HWblfAwWRh0hciF7E1ctjNlfgMK4vO3nXtKeGUg+zmm+P/dRg1v3W
K2AXRlaQ5Ulu06H/t2+KrLr0P4WifejZrSXqR99bpHXZH08s3uzV66WqDWmWafFNCbdWRv+EAcad
AhEEm3YGasLMsr2wO9jWYVo+SdWFZSC4+g+sK2g3p77kRgCnlouMkp6YHSzrTGDGqoy56CPKGzqT
BIApaA7HsJ0ayUebqiNuM0CtP4zCC/4r/e157kDiWV/VN+140of+mfsFHd1X95nogvgIinN/wTEu
VsOrqX+1wHymnGb5B1QcU2LavB/XMMkD3+jXgX9A3q53PGTZ3aHy9jri241B6g7u8NV8kX69+Chb
zF+XXYhcKXKCjgW5bE9yqAeFfTEnAWpBa8cDWPS+dYVhTcanS2icUaTC6qcLmkrAj2KGi6kGvnL4
rsd8n8lCVbTW4TRuaAiVnszYthMzRmSMTtihI9EkGBpgsClZtqgxKN2wSTQUzXN2ez0dBhlbQzpm
shjVWs8qCtCmhQn+vayNqiB+iImeM3SCsiRZdaxOzdA3h4OLxNCZTL8/LVo+8RWjOqAU4s2bpqIZ
v4xlyc4IpMJ1Kvj7lJ58yPTf6SsazsyLCPFvZ4VUadEeUBRiFH8iOwW34DosHJGZoZBC3N8KQV8s
kDSUKruMtrhNck+9YEERhblBrDFNcu9FTHupYYeM1uFQFVKIpK5fMEdBmZgZDH2WnjqtBh5dCm67
leMp25wz4sjEM8VO78I/gRZzhK10W3gIN5cr8ymDCGE1k6PkvVg9NfttMll3TtINKcVNSfJtDttO
XmjBUZ+3e+govpKCyIu9qVHjuD5m/g0ks4Q/Nu+0T++ktH8SR9nlVSHwP/QywB7+aGUCGJt4yydB
vCy1lVpfa0+/66wT3BHUjzuc3abY8gNzy6HMuB8sHeaLZRFN2eEE/Qh0zmW9mAtC9JYIthR9T1Ul
VZSF9uuzPuy9x/Kd4b3lSCsA0LhJDetOc6xDe+79ESHWA+Wc7ruaBu2T9N9HpvVr0SN7oGUUBl5x
51zoYt33cF0QU/eKuzeuAKwoN7eQVgSOBJjD8YjuVAhH8FZuVuDzu5kbtY6Qt7Jq75cyn/B4pmtV
IJfhmFj8v0MqOqaGvYa/96e/ZKN6p7HkDUIL2GyYCq+3X7UAE+VcaI8eY4Zfgsrp10vGuIcFJga6
CvYdZo7v0KHA2MC6BLGK9xtSWWQr2Axov7i+ycX3Z3iMAoPIvgm3jTtXFY20I636m98MU9ifc2G4
69TtMpTL49NBWtKUL1V7Jpxmv3epBvApLiwsqFI2JOpC+rvbey6LEv4FXhvbf4DORThVYBh+q5ct
CYFDIwrWwRv0ZdPCaO8aKsauT37CcA2o6QVKTUFmWVSrTRIx3mAr5VWdiDATDYWiIRLnK5cYbeWP
GG14lL/d7m8p0UWV/ftkcwtOTvnKiziVe+jS/rEOtJp+qF3OvvKhPbouja5h4O7YJU0Jx/JJgbdv
F4XAKJVpSgee9drFyuZ+htguH13W/hJHB5XTav860W73+DsVQrg1Hq6RIhTcFJdPD3LTL3sKnpVj
3fdKYyNNSy/tIdsJa1p7Gr4n0TAaS0oM2c5n8cPMlTb4Y0hQb80ygkn4GG7+1k7/XvidWdF5FqhI
J2vM8tKVinjpqem9x/nC4T6iPYAXF69EExcEgS7oi1Yi6uqD2eJhPEVC9IBjPJG9GJZnRqfXt2SI
2DKDGUM/MwBVI1CX3Iay1YREhYWaBrUAxprMwHAD1ehwDdc1NbRRPlOi4jsTRwjkVm2e4/FCaxyR
QiF4USc3AcLJJJHTUYYq15Dq158TUFiqUgWacTXybq/YBZ/zHyhm54Orr/djpIwJdOFJsS7Xtsf6
pKTcb0RQKAA44VXLsRw60HzioxV19ZRhE50SPU56liLmt9mqrT2B6+0mdEQufduvxuBcs2B3DaSB
C3VfPdaHeSQ3IDswLn8xsnX9MrjVum5yQ3hwtpcCJsf3z+EhER8P0z0ZlbpsxICrHqwG62ojhky2
8R16BYhc1J2ZY0a3rh4YY5veSGKJqmcTSnHqbL9YFg3RiL7N5lFYvvKHg2c9XypI2lJmG90EO830
I5aORwu+ROfVzVIMJPNU8LHMQC7UK3V+O71cB6oiY9k6zzM1e3ajCIsC2hOhtg64MefOVYkwrZcp
IBFjvhGG0Fmr0X+uq7l3yE3N+xpBIFpC/QeXr5uZ3084UnZoY5DYcbGC5Jy5I2dUFhteNMMEoSHj
9s395B5G2kVnC9QLWxiYPU3mPpt8E8mHjNsFV2Ve2Y26j/2RBahiZFMd8vAlihHBwLqm4hWWDafZ
1STFVg6OZOhxWrmFG5xQkrliPdXe9d0cm4SYdD5R54eR5EYboulLtFZSpQhxCI9qhL4qpcUyyBGb
Vg4CdN49W8O1Phxhswob5Qwcb+Q+qpM6T6pknN6c4CF/nPLY0qnwPKt6rXYlOgP/7sbscO5Zrxzl
YA6ZlO2wtfrkafswktVlBOn2me9GEr5xty0b9UHCZEo0pYhBm7+NtCOlXyOasq1PKjzHIBQAnoJu
gnlDeYkHj3hb9xYm0M0Q4yg442wfK/1DRWOEsa26qo8/jgMDCSjdohU9ujcsWMhvtimCGXXzgcIM
ICu7N96ds8nMHR3C5QPj1R7C7YT73A/DkvAAgZSQ38EinrtDSjB/kQNhwSOjLpfSFQRdV9JAdtag
5vWiW3v7LsMuyf4CBn8JO46L5W/9N4HPhnMko2Pou5nqCgOfAVxNE/l+YKGCojmF0BrvDGw9i6ep
om7mcgEjKc9Z2isBEkgdJg3cGIrHLOGJcm4QIgjqhhx8yurhURAvvfzyh6Jdp4T1wvm9mfqAwGu8
Qqgb1aBl7s9g4FCq+8MlcbRVCO6lEOkVr/KrB/O3Fa5ubOMbBTdJJzeE7VWFqK5qgLgdbDDIWgeU
TchJDWUhBH3TONzCUtD8ZMfv207cpwvI/MzGj0OTGtrPYMNzoGrEmE0/7zrQ4YjrvcYED2wg3Xg+
hexGXh/1u2F+rd3mXt3n2YMwqAqz6ObEmfB+a2hYmapCVoMNk+NKKSGLcfGIP+pvlTeciR4Ncwpd
YPwNKg/OFWK5HK+N9358Cdd1cWHjKUcqCLS+TOPABYJgmQI/n7DRu3ZCGOYGhsyGW/foHIDQIy4O
4aEU2kAydS1Gk2kFTNzSonwrQggPJVeAEj/X9HYtX51Lfw8KM7Po3njWZVWAVh1XCgHuZs5yAJsB
n/usUAAOTB26NldeUmBRPST7h0gKr1Boojjb1E71r6SdNTsQnxOiKhIEcXsR5SPHpTDEANqo3CQE
RT8Q9+gm2phxitBFGoTMX/XfRj6UxY1x2i1bDfuRKaQYt6IUwlXHolItD5+yzV98CvNZnC1LzcDx
liUVirzAwpNvXbWrJlRyz8UOEpl/OJ5/RTMvml0x+qcDwX6Nn6D7hZ/3T3bQFpBRS1DyH7kVD2N1
t1+BaID2O+BoMFZgOgnUfHifcNwIE3BWkNeQSl1RdXXKf/Wdf7cUKF4y8X6nk7KorN+UkfCgrEB+
hgvUJR70pd5Afk/9g8heQOWx2TdHvmVmBsOAFNbnFmXgkjr6mD/xNJEe9+OQh+Dbc0K+omnKLrBs
6E6nIGLUeLyApy0tdGe08Bn8mzeEiJZBOybtl4QCs3XXx9vkPn3NWyeTxJUlXKtV4N7qLYd5YKqa
wN+krEihaAoNlPXZfKJu3t2QBVPw+B8e+bTyJeaBdT3iswHSng0ovaGb13CkYSrYkDjD/zh6y9nu
XSiwa8Fma5s0fix1JY1Kic4FSN6TqucFf1GXuULPYx2k6RwxJMEt8kTUrzImQo1t7ztanK3ZzFOk
rEDXdJy7J7HWSdSSdzjHepr+p0T4AsirEVskbsFcwaAwvgyUoKxykBriup5Vg3uHerGUfkOeroGi
rZmW7euVUPslmJhEWCVQD9vz2owGmuQQvf/SJw7foo4TjKa+nSsK/vEBqDa011pEcH6OWSwCzzNg
uXjGkv5hv1s4+GHZu/7hP3xGw7T0rptr+0iH++cLLeO4Z46t8LDc9lho2Sq0ECBMD2CWEvql/BaM
wLoRNgWPgL8uPPD6zzLqdO78cKTX11+qYNe9hJCQEeKD/nKMEtUbE5q+A1TqcQ9/0Bb3fhIXBRhB
/2lQdUlwiQ8KTrquuycXj7woYwyIw3nB/o6j9ZUfzwL/6C2vRLJyAubZkGL9wqiohm1R+T3I6CJf
SzJMNl//TaEATzGU/Xiu/9Uoe6geCD2N7hMZJvN8uXeET8UsxJt/LkMse/jv+4P1IWe94K3XbwM6
Muiv2ffqMZckPpCOk99TX0AqdX+yPFipTO70/6iOP3Dg7MVaUAfdDSY6KqWr2EuFt3hAjSRgw8C0
JG8AadUKFPK7v83CjNXVDmFbn4Jh10do+jXE5lseokSgpp/VfpBuGocohDtYH5wDlOHbSg1iitb1
l6kuGcUC9/p4H9J0IjuWua3RdCoIb5W8y4agrq4REwK1n1tatLsDgctlglYcGCQJYNsSoN1pvF1J
pj9VjN1gzMEwGjfHbP/UqIDzFljpaOoXYj7Vws4G8X7UOiFHB8pah9gPmsrXQoemhxxAotEBe1dr
JHRNGIM/+r9O+qvHYI8jL7Mp2Xfe0WXwYvllUGV2Fv9qsBdtiZR2VhTS9JjhzjxME5xbMPn9dHUo
OR4xuhvHJRG6HlzKPNz9BsberZ7oqG9iys05lS/4ArvhXuQOPQQoUimonB9uYLg7KfYA2n+q93Gk
qMxpX/s2SXEp/EDPY2QWa18UtqhoQbz4Vh8ydWu1D+mzoL3PxtKAtutFo4mxtKlqQfKqEHp94fJq
S5gRgGs2AGrYVEyzX7XvTGaO6qRXS6WtpQWNnUdFmaiF4VBeUAOzL3FdviQqzHqprbT3hp9TsN5I
z/IU4xLKfIwYNcrmgh2tYa6v8PoY0kZAz7H1ZSWLWhlaI/UoIfuzRWVNdG4VQcRMu2ZRSszs7678
m4g85pGpKI0QlBZL2wnyaPimiBr3dbiUIMpa27i3e+wEobL2B+ZUs5XHpuNKI+Kk+qd3knFR6Uf3
nP79MV39FGHPSMRZVIDXab92Pwb3z2XkeU0QJ2AoEa2bUPD7E14/T0S6c7cset6tLbkOIWvf9OQx
MxXG7ief+9TFWhesLdxwyfiV5Z55+/eBe7UvQJGwk0ekOhPkxGOJMKxOqTn7YkM0WWRag5YX2Zib
8kZYIi/JtgGU/YGZw0wTg1Ehw4/aoTv9zgJ1/Mxkrc6paL+6GWoJgqu4aCYnTjocmtvQpYTSsFjp
2Ct5AibwFj7ixT00/6bTb6p8SlFK5eT3hQfvVNOvl19LHbIuuDZrBqvzJqtHgoXEQAFj+mSvDlbr
sTgXLSdRbfXCdPTTas3yAY8tJKES9cV+6XrGH3CIkJGpbWZsr6bDL51ZooVw5/r3zdhE/7WkDh1s
cGkQ++Zo+/TlTG7D5mxifPNM/Pxspt6Qo3st04mG1o2V7vJO4ahtcpZ7bH3qA89OObkFT3pP1Agj
Twozan9oUG+WQn/Bq+0DKp29wk0p0oYN7O6DtdtQEls7iHbn+8nQfY54c8cXg1xfe0tkxbQ6MCvw
BNW13Flog/jg2uMNbG0iagpGIXJS69o2jkkK4DZZ79t51VUk4bwBS2Q5d1XN2yeihhQjve02j0C6
5WL4kt1dsgTHsybitUHMdOX6psQW12dsb18lQ46IFrF6cZGSvOtgRS5Z5gf3seU0zbpi7PT7hk2p
8msm0irMIIAvrwN/GCn3Bo7yFy7C9vVAG4Mi6PjsVbwJAM7dHjFRhF6xA/hNm4H01sO5UdFMwkNS
iNBqRXBtsz9oEMgfpDF7vxUPwywLDUxE86fnQSRgfINFPswCvIpnUuzeybPJy+pO1vHA9N5LYsSi
i3E6DTZ8eE7tAsRYQBw6yn/jAHAQ/XpNSpAVN6OY7fL85Bx+RRhb2ObLjdmu0WG/KQf/U5nlJfr0
IV31Df/JdjX4c/abutolDc9bsEIGfTr8jFdWs4p/MHWSvKobO/uP/NJ9knixlWmu29yppoxEQkDA
xz5Dpzfvkh2koYqKXOINyAG7FcIZYnI78UrWoT/NOIj1dwRy2paVY1YP2vxxfi7IAYHCIAI46slf
ohRUcl23ZoDdloM/OayTlnauKQR7aHVvlKk76eLH8X5mHoXlFyBHUo2Dffg8bH6897YeqEY8c+l1
pEBI+OGDUsnLZ814USg5upf2eKoihvzPC+OhD4quPLfMLiqq1ki8FJtCCUIkKwXdUnDs58lkokhZ
JpSyXPH4Wh8DugIniZNneVGlj82Up9/ogq1q+QxLMdOPnzYAO5k8LC+CAo6Kf1OVglBbW/tmxzzQ
x6s1u+nDVNnPTTp79fF09An0bsSU+LqO0Yed3LTDA1IckILoJnMm1mDuRlMnUfaHsxswGZJxwvds
XNVJlZUSssfZrZ0kYfo0RqaA1Rs+5LuMqHjQtpQDS2jWSiFI55gOlEZAJUePKe235YkH1N3kuoRW
GEFJ9ts+DYgtk+F97k21RCSTbaCzWJOUh4+5DnDcyAJ0Y97Qez0XVr1kUiLSeEh9gEorpXH6OH7J
/fyfCEcfK9RSY4eluG+goESePtFqt3kI0P/UMnLF+Qs88EOkXJpjtwHMQuV9B9OIFlNbZRR6XC9q
y5kP+zV9IatzNzgUHMOj63pdxx81/LLFRY3ZrlxBmQ+Ibu3874GK260KtYmIZSRFdf+DU3icvddX
oLEY4jm/kRg/H/iBNjmz9yilb3qVx4n+vzO9OOHko46tzsCzIt6FMkzj204Qg9sSoQdeqRVXFNOP
8D54Fnkh7v4DBVLkEz6Xyb/Cv/MeXhew5FkchJ2lOdEHnW8lQPCw5ZIo1l80PRj7WsPfUAEVVScn
MkTNEEpfRRT1FR2GRhd0PrMnrV7+PdLPMaRV8815No9QhySK1T784zyRaaoTKgatW+naMYCcc/PO
y7Q/RZZLMzuThn+AN+AAXwevNRkLalInpyQM6SoGVGkJrB0yQRkX2Pn92P4KLJLKXKEpmR/VOpxr
2p8h1RWvs0lhlPYcSjdPzN/NBrS3iRhSBwiQF+F/jWoZHL8FhwH4rDMaG/rCrKpwhd997qRlX61g
CF4583K5eZSj4sTfX0Drg3+//9tYiry3xKXt4OI+C2l0op8OOHKRQJVQLqq77LweSCIt4IyHlySb
jxSUliAe3VcfzTUtGU7dGkf9AZ1nZvq9qcAJ7EDFFDeEw56pVUOrLKFQFpeUaZHKn+Char5k2PC/
LLDr3LGWGnxevJU/14PDwuOWKYwFr2zZzJaYgUoqwUechWYNYvtl0izwhT+gsWUPkkY8K+mNv8x1
kKfQ5uhtRpp0tTaf8rN4FvqGB3Umqd3pV3/mzuznGU1auTbpf2QLtxL+LCT4oW+GgNCzOZGDp8Ge
HnqijxDNY2VrC3UE0M+CXh/yGbFrBmbvg4myjr4vClIvv4K5qnQsvL+kvacB+PnluU1eUS6WsBJ1
70MrPW1zINbfcDG99TLN4XuK2cICyzmYbYEfadrVAZj4b3aFhP91gshQD+RqHFfqBy8hOd5tg39B
6Oy/Rv5aqToT7SWPlKCxhBrQUHaWl7DyPzl/BPYcuoz2/ZLe8AYdnj5jqbdjLRmdZmBmvmKoN/82
izz3GbqF5KNNe9GFmXUzggRXjK210QaikQu67qWYT6493hl+kWnCnY+DX5znZYdWDeMGAz6/EDGh
zjKe6l49a35+OqmXOsDRxPHkRrfr8iC+c+7Pc13Tnxu555FY3vipKcBJpeHV2ObB5PAvdhrsCa0L
vdJZK7eFV0u5f7xs1t3pyuVMaJAUWYVl+v9Pjd3sTx7y5wPtMLu45uA9SeMatBwDSBhkAwxNHpdO
vQisgHk7lDs9jAotC2plWrnZoiv3Mn0HIiqiqQvWWpJ7g76QusZIbSWHPkPSk2c3Itr22TEUYQRV
CHckvNV8685tYCJhDqDK1MUvGbytnz0tbbXNNvKCIpnUEvKsOCmB9YD/g73O9+V0W1MCCbokw/Ok
1qHh7qWYcxxOeEPjyWP3J8fBu/HhzsLWMhPoK2D3jgAM06tZP7aNxKw47GitAqCFgYkzBNW9iYR6
mgzsQs6XBXntDQItScUDGiDI2Jp1CSR/kJeRgbXPpi9q4zusUVR6U6GCotVgAYv+gXNqRFb3zrGA
yaoCvSN6z5XgGSBFEaE2zRe1Wan7dV54kT6xQRUMC9ATDLsb35wumR362jkvSBJVsjx9vORe1jFu
Se4R4oT8jTNJDXH3FWO2aJHyn2Eo6ONr8wi9eRckA1P7LBbTa5U/W6cog2jHubexbmpqptdxLgMi
WeEsCLuYsDex2f1hYMIiajj7IOiIe/6/sa2cp5xXPhWN7wa2QuaEzu3lgQv1BVfGe5JA3AK+RnAx
w871LFcdplVekTYGek3j2ODTpNZ4Oc68zgq6qwvcfQr5bJiquW+cssMdENozqfj0YjRU8RHYX3cn
slSetbH6PPItM0c35mnAUbuX89vQFPG2F9k0WSmM5tjhHYDlMts8+cFex5t1VlKEhj5V85vkUPKv
YO+Iw7MasUnx3RxuNeSFg+T7DCDsfoNMqGbQcvV6FzmLiQ7VCB2sFHI91O1+ncv8t54EcaYGW8jp
9Jy8lLJFq0PdfyEvCc4aYgNJFtej29nCZ/Nc0hJg2nvf9U0xFSxEG4P0GfqQXKKBR41TvdoIM2rx
4FkBSDyvXXkXiEYRCz7mMUie6pYCdUAdqCZfDDgtrRufvw/zEtBeL0Kq7h40sshBvC/oPIEaO1PS
r5zheKmfwHxnL2YKXSpFXV9/IriruItQWdOufcUiurB38UdWFq4mraBtFBGiaRYx64Iqk+PW7xbX
a7nq73/37Qd8kQcmiWUaI7tRQws7o9gnpEbWPVVqecvW5g7mjmvoyEOVEglHD5NM26x+Jt+ED6ku
2vzar/s5y/CzkkA7bzR4NN3rdzdxiWA9bkINkTOSvgtKvakGRoRO6pHnjjSDUMXb3EmVFRL1cE/1
XBNR6vD+Y4AbA6UahWb1tpVqt+D8D/ztn5c+r0WReS8eQTvqHKPhTH2KkhF2xiIXsA1WMNy1U2kI
XkmlvHw/W5lOHHPiHAtiyozm6NCxsPz/n2DEOBm3YPKqC01bSeoLBUo3uG6LZjRWG9UZ4dg27TmH
NJS4IafLO7TpUYmLo20FZsqw7z8L/3jekNbosS8GwQfymgPqryl47BUMev/IJ6fdw+cdvhoEYflq
f1Irw0+JjDfAVzwAonBhvOtEMoYOMaldCNI2S9WcNzfSTm5StgNd7TDIMjoDym8xB7uODidYvg/u
AtRPsuAu4nrblbKp3iGGb+meGesr520NZNSwJwDjkA/zLAIHx0keRJ31U6FFuVRc7Slz42Jm+aXe
N/zRDof8T68gxxfBhKmyZTR7MwnNozCYM6Dpzi82E4urNt28hopJ9ez/QIFVDpaxL10cQ3Cg4HsH
SVgAYYsCYiYKmwyTZtcmG94c5esYA2FMBMCGm9uU8rIsT509+tfVoPvIrMTrlIIJ51QtEzg6CQqf
Mg0kp2R1+wvCNT5c0F2Krbr18yhK1+3pL950dfYQWIU7iQC0Sbyx3KQQF45w0pH4w3CRzR+trYz3
X+wGJQ3wGHuJDFPCrs8nLTHBOROkxFX/sjAgitybzmar/9mCOBFU+/v0P++WHzjADY34ZwQSaI9M
PvUVIUCY1rr19s+1/Y/sk8twahH7UtTl5svCrmzZdJwoCPZymnLEfRNXZ/0w9tWjSgCohnFW5A0y
6lmIb3GX+63RNsfGYtwDwhnm+CwQF6N5Pl5u0J58BPpyBarFaKvhBYPcw2y8WqtAFG8SqircHsWG
3u83H1jvUFz4ue8QTIzRql03H4ynvTiAKMsLMdd2XE+B5lOxf5YLe3TzpxW95Zfcfn62dk7Tybf5
b5OewdcNIwi1HIBhkFbcNqi1Dw3UlpQx9W8+8Z25pler+Oyd8v0kxLXuJMrAOFR7KpTs3Z5o4SS1
w5SEHOf8B7LJcpvKBuBBJqxA63uhKfcjyaFmQuxuzbfmi6OR4xXBoy5xAuaO6u8gG6IWIKbZ/GgH
eoUgnc1DOPCtP8l8FHhPRo6QB6ieEHpYShUL+QWGCdDKcCfX6LA58DOEQjwsqah69Ts71jjrxda8
zzSljsogIG5gI32PQ1S5/CVz0bW2aNzsfMFgN6cNofjSNdoBRVaNoA9fpTVRNe4tOjvFUSrbnVmv
ZShf1bBrP59wjXDYfxSHfd5OjCgBj8t2dB+HZfOsnZMLwJT4XF2yqPtbS6iInaaRybY3b9DyWM+K
IyTDMhmjDAs59M7OpV2TyWuLYxByVNLeYWF60B5E/O1wg9WxADfiz09pzbCPtXCrIfdHvlgxTITT
SGYDUJwj/tYrAT9hP78IWk/2JKCMfV3XXavtwKJyZ7pa/08tFR5w3CojxYbbnobK4Ref1dccFsss
iu8b+JhczWfSfnV4fQdmhYeaWu8BjmJKaH7tQnu8kM6gxHMYhcB035098zJHmJladCjTf0ROZrsZ
p3VjnKdNZCH5bkhHi4cfZ8Ex8Qj6Hz+VlDDKQxDq5LxtxWnhET4LGp00ykczrFqA4yPlFcRs/7uc
LwyxirT5M6mFn77PRrntfDTCdXNeN62VCY+OLpjV/7DYtPwazX/dbMxQPo2lOuXDCMfyGqz9jXvO
6LuiPKnKzub3gJNFhVKxb+C+OrNHBuU5m7a0wBY70W7vgrw/iVtIc9oDZ4Nj/63GetxKjtpRVDbS
klSSRvnFjOPnbK/k5xOLVN5trPZB/hcRaOtkHq+mbABNsnalBI8ZB5OWtp7VybxJtBXbaucLAeyz
gASIzJ1mrkiJBgqvXeimtQfg0o3YSxDLW/cpv/LaBcyEEmf32NEhdt1kcK9pvhO0fPvnq8d64JWF
atjBZmrxQbWM+10EKURWa/4/Jcpcy8xhZhDX0LO5MpsgEwTmC8wrJr78Sv5sbiK+OYhyZ9zGE9ma
o9Y7QATWOZ/nmJzC1E+BNJrI4qlOzz84/5lWKqMEiPxBH6VhY7QXDmPUfd/kEwtFFftNu/FNEXR4
Kdc0G9oYjZ1qqehZsqC9WiPGP0LYk6h6jA250LGJ19Fqmx9xrKdN601mvJqkBK5biMMVYK4WGZYA
9Bafd9YIF/Tlqe1eelOSHN+0RzllibaqFRwiLyTZ4uEwdBQur6PbkJv45yDKBkHJC7+pG8npnW4X
4zsNXqMvB/pHMnZ5mzORwaa4E9hFra5MyZ3rstvLuLJGnxkJ4hJpgbxHL4VaKgIhLycnYRBIqIau
JxG8MpayfPQheHWQM0x8L9SfzI+OWXL5xDfGwTqvoVcEQGjgMeTw8pk+DWcxhbwDrWnmbzV2QMUt
RD4Ih5+n0qgF/pV3iUKalJq1Xfnj7m/WIIfKkONMpXqN3RKhKt8SVSLaD7ei/QIVOJNTsyr7AZYc
bWXG47VtoW4LX8RT5agQQEpU0dEH0Cg1AcHYT2GhRoAtnVCge751J8pOvvNJRcXNuiAoM6uS8wj/
eMBDiJIThr+KhEo74Lg+Lbud9+W/noZD9S2U5jK2/v6OA6/NWjl1snJ5DTHY7Mnh1hRXaYwXDB5i
0jBSuKv+Xp4ZUyIrbQJuvvZ0IcUQP/M4p/NdCJFAhvie9hhENR22DgiUfyANvCSP7E2ciZDRzc1o
SIEtQJUSgsa53Ysmpdz+xfSX98hVB5jrT5N9UrZRvvkwr5txUdxUMTxEPPUtT5prpjtxRhzwFbbI
ECkJjdwmUk/tg6ez7l+94phliqro5dtX9qJCUO7BfauYppWutVyvQhEjfDRoUp+LQGgkN94DooVf
xpb+r746KwnSZaQHsDifOTGLdKrX7w9AQv6jvqEBKjtmvKLJ4UAnfZqSa7vJ5KH7zZuDuGqP3Y/I
foncMxCOO360Xgia1zVzqHaKAD50vlyOEM/hHOLUue9RIC6WUjmuprC8/2PzE8KHqWGubkKlaXk6
XC2O+ycLACwnjLaiGEUaRKwo7UKFvXrtjU/Bw7ZKhOIiTrh+4qNV8PhIbBsDEaob6SRbl4+xVAJF
z749QPjljjBpktVzDXK7Jts3TflAWfkPS4AzAonKkvAweF54lY5Du3DX86Z5lfqqiu6poXVceZVJ
u7CJelYz+4mYr457yiVLZB+yjmRhqjGOQUzl5+kIrmj2zA0czgVg86LCSrWH0/IZNUqFsq/omhoU
YOrD3d89fmgf3sJtXKkEL8UuMuMAwapFE7XLkHDkoI48usAC+mCYMqjecutFsF1AQ8E06SasfJq0
N+TilqVTkICFulCc0DNJ4tCs2bKw+yNCTrA9PAYd+2+yMzu5G/uWv8SsQfHBGojeuawcIkhopHcd
Y7eujzLW4Z9qe9o8v9KCT4Bibr+hDZHZ7hZ/EvjtN2CNkvwM6MknX8o3rX045KuS1n5CO7fl9yVU
+6SE4ilJ3kf3uxweLI/j1I/bmHYsZaxF6b0217ftfYqzRzhbgA74e4iH98VsuFiWBmVCvy/+RQxr
Vrmiuy7pkXG+QuHWvk0Rrirol/HuoEYSLU3BIccOUmWbaaQrF7qM/oI4q2OoNP0lmOUB7YROrHW7
qoW/xDeixh58fdeliQrXkX6zppey19TrWYl1sODDHYxwF+58GhFxZhUwwpZcWC5YGG6AzNk3LXbb
Yo/uS05sDSrV929kcpRToVQmBGaXah6eOY33+y7kCvvYpQyikmooR+2NOiqA94Z4KGX61rJtuAC1
P8zvF7LJ58FNxFQwUoLGlrb9m2g+z1LS4jiyPJCHg/dxf/2ZtKcod+DAFt51Owjsv8CF8n1/NIOU
J2BrAL+6qrfpHq6aUPQJtaPJpO4DuPNDLDmDx4NfKR09g0v6PnXVYFjQvjYcX+DczPSTu/eUUSFe
W1NSFJQR5tckjfzIHS9L6dA7IUGaUydYTIiQ7jDtBni6VzXAHnZQeAfGbxhlOWvxKvF4/9u+ROpa
dkuydPykrPBOFsQ58DrKZSIKm8+yRDS38pLzw38F9ik2uVYBbW05wp/kIGYp9BZTn+5Qy+JW6xJF
zS0Mow9huIKsTLld5LukXxm26tZ7wZMTYydLLDjI5KxnBNrIApIEWIy5gXsINSuGRttwYC65cqiV
cEDXuAqTTbbJk4naX/vXZnalSRbgDT1WbnJbdDy0oeDcUcgWWM7Vn+l41NFO1By3Wevr0DC4NkDV
nH88Lq+gt+03SwYV8QR85dcTPFzCVeye2fdgGGHcCSndal+sb19x1qXL4WHBfmLC/2mZLHr0gZR0
TSoYdr5eA6GmXwQQZ79Tnfjrqidh0NkRIRn7yGY+FMh1Sqa1FyytO0o95HAVCEDCo3aSsXavTQ64
AC0owH1Z3xCd02g0tNyQQQLpl3Pe7XenuB0H661VIas/tts75MVBapy2xDE+TU1iUv6VeTMs6zLL
KFFR+h8GDYnHMbn+pKj+rbeKgEWElRntpU8mb0n8l1/3LJwyAtIHF34ke+NuKCJX3VsxqdsWRCth
SQDLgVcfwUPzf80TvbLSrTkvSEx2hQ1+S8ZHq3y0stgDzoRr4ikERRoqDwzSgW0bjvr8xggyaUXu
aa9HYAgxxWVUN9fbA/+DZtBCFgMwTAxsHGtgrcHUKQxlUm8HWo3O+UWrkBw5uAUnL4Jgr/vORhpu
0Hi1lteiuJSdAZ7TQ1GH77cf54p8wJ3RZ61o9Ny6h3MBOcEeJBnQIbOehia3d540s4QNhyKwDjjT
pV9SuQ+k2fAeZfYRZ1FbF7sO3UN1qa6dwlYUGUoxjqYBGMXAZu0vJ5mg9gqkVwBPPWOxhEhsp5NV
ppBNvlyG5TjBAzXY+1zQQaQQquOgbGGb7JYkT9xsdyiEBmFDVVQI3apJ1hETQkgKW+B2v2pbXgHf
TaCR9H2TQcbUT6Q39N8pNlYIC6Lz3JGuG8Ch/YqXtrrVXG/h0khAaIF2npem6RPI8yVsBi8ex9cT
l4LJC4DXQJd/OZBljyx5dsNcaBvS3nP99f7xIoUVDEPUo+1/KJiMQvtyEWGnvQbwVrvEIRtFef6C
Ea9kkXgJuzSofdbAezLzMwLSDvdyMuZhpKx/cYpI7IJXOx95opT1Vs43tuq5p4vXu9Uqv1WGudlQ
xNqKbWPfIl6JkQ5xldm6nPNdQrUn+5ZNLkk+URjLpvMHew2od4nD6laMRzxKGpGlTqr+TlXP+Jxd
Rc6Rgs6ePfpgRmAn+8G6Zih2oBVxHRqqr5R59/ttw2YLbptAn7pgrMbcIFH3pxRZ+b+yLPnP1kCx
rYhtuVrr8KNge/VabGdSfNEub/8hUD9ttPomVaCotafL7wDgEHnwN+Adc7qfL+2DPfCEy1iqx2H5
763JwHlHGDpJNxaqhWRj5ffrZesBRX9AwBaSP5pYEQqk7Kn7qHLVnhEWOozmo2chb2r+IutKt8xC
+SHC+DXJ8UVqd/9gUokh2o9NJg/2JHSLiRtXUNpN/i87VQyH1lK4p+a9GRW6PR9CagM5FcMFoVkw
+UjwSuBXNRO/QazTX9TzlgO88b+N2B6C4xa7cEgKzVQn/wLHn8RPvqKqEpNU8SHX+GTB4H2t5bcM
u3AHAiYbE70pkA8T38DjtRzZGcj5RtoThb1+HUGSrDWDE+xNO14BjI06edX97WQ57BqNfOEw4o2t
/lOSxkIsMPXwNwt2nwbHClMSKp3AyKqnjElNJeNoU7XECicl+tm/gNi2EoDpOmBfH1zJY5pMNwOl
xYypaghamVU04+HsVO8geH24Udze8cIjM1V5ZxyvuiuOBMC2Twp2tkG8755GCGYro6Pcf6j9NKjg
YSQjMeqDoeXDRkkOMs5oLMIABWndmDIzey5OhGfzIp7VaFgmZ0Kb8z0d8ugg2wNxL6I6UDw4rXtr
yAIppTEvn7oWyHix4pIeHiJCA5FR6pYTY8iLfGmDoX8ZaQmn7fZzfZv9UHIJahVE/ey68HJrxO2p
NHrqIwiIWumEgCjNfPeOLI9ykEsUwEDY7f8wtpgo2inNkLZWMBHg9hRxJ8CJrUtFKhBBJ0PQ67qf
1p4fplsmLRUuaV2RtW+n+4kFT0mNV5Qs0yWEUepByZz74cQ/srlFUgZp1NyirK5vSkEOWbUSaITx
7jPWGcMFtqxdoW2+ZIaONb+jk2AXTKJsWmUrwnah3YCcf2KVAjTSyWXqBrdQ6rYbYOXnidXZqnD6
4cGP070eltc1ywrDM43WC2xR+gMSssT5KYnBIYv3MgDVM+Y5GSRaIIIPtXeSSJn5zmQrm7RkTlr4
Ut8R+PMRuoLWIR8GqXBinXgxAwnLN+8BN348CKhJHdXgIAgZWdqmLJ+ZKrN6+4p7Q1Bsx1lnXBcZ
1Q3JwQK3rB1uU/8WAPlR5aNuCBfISSmEunbQXmIuiMaQfdlbpk5LL5o3ehs0/fpAwAECmXUCIGaG
ijXdNRgEPPFBAPR01w6h4hu2s87711xDElQAtYkwMCNYP0ffStfZVQIQrdUTKOiuhmeaz6toH52z
Q5syeT//hcPUhYcPhurUt57IJUEI/d5w4i5CpyFPSScfoeujMVYJXk/KkU8wAoaBhnY7W1vdJIPb
dpb4DfexkEOBBFCxvAdtK2+1YE3u9mYfOS42jaDQwn5ghubSYCENTJEMY07WKJHvwGjJqoJWUi32
xA/n41kViHBe/bt8TKnj/OnBeZIAgPZVXUQvAgdG+Gt5nPOAtIib8BhgvsWnXL5nnz0WbBeke3n3
9FTvr4Am+2b0aXcLyI7OyIq+02J8LHVGwLfzy4dpn1KmAqK73PggighAU7jXuLOPV4vf6HqWBECZ
Afc4Xa4/MHLw5STy4RlCvJ8ZgqPbyKejkygVDMFMPoubMJKHRmgTu8m3fHU9XSu9ob5SvKLXAcnf
UHo8K3iANAgKqNJHmlrtc5a4GRpIbDv3aduUvKVg3qQ5NsW6awptVsmm0kUpSk36Ov4RLjlTWdVm
N1o8VLgF2WDeCJ7HYu7ZcDC51bqdpz7jidGAsWEvWY1lZdTgRLHo834fOtNe+uL4tE8pS8gRXeg1
vxYTjA4X3nPawRDaBfr/82tQ4Msqjz8WHWulGSiEAbkgdktiQobLQTGlRZKy+YbpGYn7SnNehC2Z
cf60biFVj+hHm0Uq2nFtV4j5I48KS3FaR72HU3u41kjsrlEeVP8pZ9XuIeTHaCqtbNk0ZZrx7HWt
sv8+J0KZwblSLqHgO6MOaAEo/4+vrZDeN2FVRhQt3so/xIebmzRnjEMzPJfCUFrRFJc1hYAbmXQs
dRguXW02G5MbnV3rGQkSfUiW6ycFFY+oIpTCbsdVreclDmBrMHXCSDbqlFJqhcj4hyZVwB0kQpyb
CyyQa7bKpAccl5fVovWuK7345ltgSIL81shWDX8X5PzqQZX86ukelIPDsxGsK1dGp9vAOjo2sU2b
AYIz5s7/TjLHdFci1ouguC01bWWHlWew5dBJwquPew5kckRAXuDJTIYukajyxLp62ayb2wYoFjVR
9JP+5QqzacMaKb1O6s7Rp/5b8sx1RqaJY0JNcDfSrAm0Dh9cbnUPFysa0pf4SXLK2JmJLPz4uboD
yVpL20whl0r1xWb9JOW9ZEjWPvxDx6pVd9DpmPIG22ProRGNnUTJGsLy6I9WTD51j72nojnNN7Ao
T2il6+DILOYCGL5+oQHkfru8f8EJeLtaE3Tm3ynB5PrR6ewcJ4gASzsML9ya/QzW9UnSjl6zvUq/
hF7EWTC+aJ/t1vNYD27vOq3bZc+wRDSGLF6vBkrTuLmHL6K2NytRqEKQeq4r70CtzPNJRPEkaJoL
87FCz9TnlRosT9Ei7PibyXxzjdXMwmFj7CkIV8hfcOaVSYeRxzqTveZ0xG70cs7ZCyrm7aehEo5u
CSfGHB3uwNS7DJUv5gyAGintmn21kCj0izgtewl7xWdwRLVX8Q4LWWodyujJAjn5XQoOnckEaimR
NgJhcH1NovknIUKzeh5mT0DERlgEA6WsGhw1MQCtgWezDq9Aoa/BIOwP1rLsdTKcYILV35Q+TdNu
1ruK5cg3SWtXncO20FAVcXRjwOc6ndLMmvu00qTx4KSWtf9thExpTRTiG1ItvS+x6U9jJiNCmTjG
TMqZed5NZEE2H9emXUOl6GUKexhna4CkhMzeW8RwKjwqsEnIseNWexQVD3lIkxUsI1jdYC5MkwBW
dElL3H9ayBqPaRGdxeojwRNvOQ1jfo2wlQHct4lBtIlP+jWN/2FeergLjs5SondI/CzggGsKCWrE
6HaV8sA8fBzlbcgtdr73CfANHn2fNjvYObqrOowShFWc/ejXTm6nVepX2/+QWldzyWEXcLV0TA4o
lglZFKhRz4/wHwurS6C8bfeeo2ukIZcd/BH0MoMKu/wZPnjzYmt0Uf4X9MfegltZKfsx6apEPvXM
HLlAzs+aOZJpEVqyuEAbH4M9KNvjgWB8v3agTBVR5QpF7NJ5+vxWBL+gKE86g6KgHczxVyVUb6Qd
VM74vsFdweXA4cTNaEcPf7N82dCwuXdDMFGS8FFgtmrzJCLI2GmMcAVTYjG6IzkeJSDXjhwxGkWe
EbzLGb239cQBgqRcDokBk4KfFPWdjzbWP6uHX5pI2L/Xd7iOe/Zs1ybn6un5Oz2ziBA7VVsZwma7
WTLKf9ikMe426jNiRnXJ7cZIC1Q4cnNgut1mdWrJuzchQPm8Bo2mFG8Ng4CdCKT1G8ZDakQWlFJg
wpdu7RJjF7wt1w3Yvd0viAbkTsb+1tCe2ekh8UJ0gCMGqRuC930w9vohVEI6l7i50Xtk6lDMe2A2
4Tgr7dZfoQ/xuW0n+h+hSnNYEN0VLxenv/XAipIeJSo9Dk7/wNNG60LcinP4KwO0kJQc+etgV+eF
KKV3fUCSCX++JhpRyphNdv9wRSvdU8dWPQFsgOEgeAPxDFNufg496XYv6eDmvIfG6LtQa1r9ZaoM
i3QNsAsgkwlHulH3UKaEGcBfKydSMUWCiFXxAhqInvNymFojWQ4NRMQKXEh35/1sqQILGcWbQ+DR
Ypj36HofZC/dy1XQzN9Ro9TVztKmFbHMP1AGWCv2lxYA/P/EXqtCQ0Ip//ewwhv0Fk/sH/A5ujmG
Md1udEMqkUHDZVyki2g9ToLztddSRMMeociRlcStUXA0X0r7MpE3XUeDEo8wcAaJgA34t7KdQzV1
rjizTyz+9ri9D4ll5xPRoPs+TpeU+bDLtcFN0qHv85CG0NKcf4nznDCFaRufeLLACB57Wswjpr6H
K0WhtP/YuGzEpW/qcYCTj7uZqbgBfD9wNasZMILmZdGEmwSMD1fcw/Ug+5sMqOhO/mrpAWAV0lqi
35psiXG2nMdowTBKkyI9QR2S2ptVAWtvWK0cp8jOT8kTAFMfZNl2+74wNoQDQXDp+ZM46Q49O+U1
9J4QrC6xRQwqLG3kkrDd3hfw+33llEdcLS1JHLwm2Wki8XtNquY4QvOjNHobCkorTQlmjLOdzgJk
ad0q6Gs7DZeP5DBmkqUOnUNymB9BrprblSqS57UXR+qT5gMdDLxwamu7McJbXxOe+Q/bchTkOy0w
8NGnPF7qmTB9BuTy5SWYwspGHOeKepbZNsszcOP77J+qIWpLl1ePEDtZeUe69pl9jIziqClYIvMt
XeLAtAql6cga+h3DEpMwhXdRolSUACW35zoQME1VcMuOg660tyHpQ2tjIVCuoW6a85o2Akjnr105
SkVAIna6SDT3EWXMRrJxjsgOWjJuu5mNP8WG6Uw1zixP4J+0HRBsV4jxOz49NSpyFnSkAhrNOvSl
XNDgpVuRoD8qU5I+XkHordReIOo2wcvMt30w/lglZhAAM1HnSHmGyGsVTAH9zs/ImsqILPNZxMFG
0VZ4i5KD9GnB8kNuqfK+pBlgHji5udNO7+Vg294uJjp+KWNMN9vsjA/oXAKK+NfkfjcFQ9QdjsKn
YNdC/YSnMta9pYDVkyoy2QM7ZBjxZt/XFeflYOsNEmtkoBJngod1mj4rugffDCVfy01s1cfF5FrT
lWyvTSNvRMzVkZ8B+iYLYmAEqCx6kr6ja1ILQ6f3blALyAZKAas6pOELffO5yPmqTVottc4im5A6
bX9/KrQD/fUBVXxjbTxKnF54aGM+seQYA/28mbabeKUYG9Yz5PZg0uREjmRATG+6XdanILNqs5Wb
PTNAVe9qnihiiNONqzSDfOsgkYbQR7wNSk3YXTKvfrQHt3KUbs/x+Zy1dWzvH8Zwyd+3GgU12iD8
y2PKCjwKSt0l/6IPJDWS8R5qGkoOEg/nrMo1/kYixmM5QbrPy5chzWcfo5VEECUaIQKN7y3ijezC
63DC5fo0CB7PJOkadoJrq/3FdVLmvY+Ays2JVEvh2rEsicYKSdN+TeFiFdVpvIF8n8+xXSGTA253
JecMpgaNBx/ihDGqAcZZLMYxPr6IbSwmUsGg5vootxjxjv5kwcSu1EvI8yzDKvXPRT23tKWCt6iU
simw/jkmx1izdk8oU2VF8OohT+s4n2UXlgO0PdCveMskZ4IJo6mxzvQwtLaAz1msN9UO30TOpcaN
csgt9+4lT1NtznFstCzmA/V9HHXsdtBnXmtkIDar4pd7rDOvHD1hz1BcydZNr1HYTJr6CLNWb7UP
MPG8QQ0fKFumLPtfcwFa/qBVrznRbeLzVWUlNmGSm3FFpTz24ialrJtC6/lMK9R/7YC1V0bcL43x
wdsx2lq3Vg9c/2xw9jmLW9z2RFJfvifu0XjxCsaKtpeWakQXvVbEpkv9G8NFjsBSg3OmZl6ZGKx/
GdW8FHix2R5PZtrUp27s4jnEARvqebhYyq4gwEr68dg9lcT4kiyscOZu5VlBfoTe4HkYDpi1kp+o
g0qHY7MSSLVjI4wbQO2FV00oOn7kBAiqSZjEfaxKWap2Wj63fJSh1HRDkGlAclY9tPp7h2MWadiX
IgiykAuqaqPpD+0cWsQVAtTHnritaG1uKwoK8x4fiRSTq7kgAaIUl9Dt8ti1PH2rhlQs+/2eRb9r
RgTqyzAkKcofBw5WOpb7fnIswi51LCvbYYUfx1m9dCqwh7scxi4/qej2YnZsWionumpeLxxdFOUU
3jAE0tE9yveUMCN7G0OEHWnD6n46ukDjGeTpTIr6uhVer5O+srPp6860Kff1XgXz1VZY88aXpaXv
cGk7bYEMv8U4ksa/TN5G7hpTQSqw+p/Bu3OpyzrVqFq/FjvjrtIpf9CBSQyKHQ85yVxOoBtiRjSk
CO2Sq5kywgVqrJrVOTYzoMIlSLsDATztf9PtZzLGxEXxJ6fGhzaELatq1ewxgZU6Wh1JxdNF+tJt
/yE36iu7UYeCmiJRrq4sx8Eel+lyLSseuBBPu1g6lPeRlX+0KMH69LVhVyCWh0ylLsRsUbNYvOl2
6Bs4vIDkF3+E690Rpw3xU6GSkk9TojPsQ/xCNrhgUzmsZEbAlev2S5KglFFNjYAc3F7JE4bPgg/i
4tiouoyRJJHrgYr0mj7ESjAVtzsyBGqaxD/1PGhxs7E1/dJGhuUw4tkoT3Us1ylLSABcmRTSWTsK
mbXjN+WkObknoXkGgDvckfaqI6SC3CDQFAI8uRn0SJwaAQaVO8Wud4EWyyBVmuSxSJWYzqHyFPpw
nXSzUshBV+4g8UZefzGW68dtPHRQPwGbRmaLZXhVkoLoHOCYGjCXdffgQh3Z7A8cU90ULjP4sow5
ZQr5UBMjieCJAmlyzCrzkunlmp3X+h79SraJaIi60wf8wk9ULYXYfM+MnUcFDI+EVKF0P4aens1E
PJrkzmdmJ+Cd4HxL8ccYBbM5LTzs8KE+xcEBQZ//91+gg6k47HHwRifofo1M6fhl4urrR/yoxp2B
RvShrbnRnw0mh0y14R7K5+wJR9VvpJMnVYBPoMszrgoOpXPnDw9KWT839Nl9e3JxkzpwoUqsQ5hM
lDTLvOWdL4/oo3FQ9pJiISH5WzvH8UFjWGsw+h64D47IoSUSyA3LmzwiUBRbJanyC4GtBgwbIk6R
9wwBBP+cTIkeFMvcOVH6D2jCA4bHfTT0JUKABt5yN+1aREM23Feh07qNg39J2m2iGPAKN432/GZA
MRqGmT5nsOiS+/HpuBrjYcUqsR4i0d+/QqjYtkHCocQULPo/ke7IlYPAbxB0LC39L1cdzI/vUso+
eSizxbkEdKU47duMuLL60woUAvoJ1tMBR1kni8VrIlxIHke/oXAOUk3dohdOPVrDzoZPMqqJzS9q
VjPpycmH92MGwhDVgSjvju+VIw1JDT/wL4oE0eDy80gg8na9tddVIRy1PnDkHa86el5YVDGg936Z
ZWJB0jDVqz68/IXXRHR3Gg9fNpEr09X6j5OwWppoQ79vwpmxovlrmsXrHb/ycZdGh0fUmV4RK3Kk
uQKsuylP4wmQRL977ZocMy9FwIizneRaYRC4X5VIQYBkS0mx35LVbbqlML0tN0Era6nNdvGM1q8U
1mogTtnSBp1DIBbWZq2f4+RsKUPUpy0IlovKndE9fTK88ZWW30vDqTwJV2kj3I23vJ6+Y1qnScM+
S9I3C0BHuinbnVG/a68ZUqmYTCdyFJLfNZ3vOTU7FiswkShpkvrEud4APCIUNyFQOX0tMAMPYozK
a2dNMd3lcRHGRFpnGrKdSgAkAiQtr3i+YsmOGfF7Ww4RdkCiFvyJqaKCVsFHBMTq6fGi5aD/IxZU
JjF35Vqy9fwA3AaecMIJXDXaWmhtJowMcFfm/VfeXc3i7W4rico9bkxg6GBRH2QKWqt8T7+jOuIb
V7TQCQa0gjcJVC0FyVmnCNSdTDK7xEFDi/I1nvgWuoUtAV0zUVtWqN9IDZUelu6MsR0/IBMgUqCs
wRu2FaPPoteXNaIYMR9OcKF6p7NmQykwO6nyqagMCsQM1hw2GRsB+12SyMXCCiAaYFZlMKuK0v4X
ZVFYAalaNiBKbmqjCMU/+ZwR02b1AWpw/ozhS4HNR3sX9Yjp5e8BtLI0Td7jarqgyK/4DAIVQ1jv
nv3/iLIrTHYqWqstPrQy4MSBZQ+tFSRNXg7MpNYkib3x74LSoccPGM3lvcgfJyF7yVRHL/4r2kP7
irMp61S3+FAYm9XwRbsxdPnzcW8RLawJPsZBUMpZqx3TLSzOm48713+yD44JhiElGJoB+AYN2xVX
KjbsxouBCp3s/7grYxnDuZfHaarNGS8DqwuJc5Vx62O6OeBLy8nCy2hD975AS63KH+sjiu5xk9SM
5ycj5y+q6xLd223XzBoG1EDdMczeKkkDcKkG5Gnek04VemvW3Mp0NFIGOvAK9xd5pma2dPsOi0mg
BBCvY3YUvQovOPFrJsk9w0KIaaKHrPn5rk+HqPC5NoSZsm42IavtpglQ92ZncYMV2jR7ik1TIJlx
k+wTroQpO4Lp4YZ7gRw4VwE1xv59DT4v/kY6AjUXoINe3sMfOdi6bBljhKjZuBzseuvi9BSUETpx
bcuQUkkFq6jO3DhYOjCXYPP5KxnWbQjT9Tl2x0OmHwDSE249/3/wuZM8t3dsJInZDb6CKVLvXLLq
E6DOMRw5hgoz7AQ3y17Lls1vHB067Bv9Qi1criLOpVz3sIgf0dxPMeyTN9iUlkeCTvpTlC2U1Fx6
P/1u8CVxBFHK+RbKYRuGho87Cr5E/tke/ZtLC3M0ru9afuJTumfUWFK78kJvIzWLmlChVYK+9AKI
FOpBkkOF3nVKClz2x6q+tqBeEqCgLmLz7UDveF+GR2+FVbxE7PauPT9aRg8s0jeSXUeeZ6UIy59W
/VhmDmCVWbq58OdYnCdsRHOYobquVLafuRQPjlWCbHnSbfXmkQAw98YmzK8Odb63eUZyN4s2pxSb
R4rblaZHmgJk8pY1sgg8iZUT/mMQlOCFJklV5sBMlyK/Uip1tOyFB7nF6TFmL4cByimf55G96Wic
7ybt28sxhGpuBWLlfVs42dKtQFa8QvnltJvWGAwXDR/Hw/gzE/esFhsQXFtG/MAN1Lb1LCpqUgJF
OWDhxW424HM2Uk3aTaA01xqOZmRGZPniqdd1t4JnhQs7Hcg7B9uV/8X4Zsk1R14/7+CZwdGuBQ+6
U8C5h8JDoXFNCCxSvnlDtkAH4fNIiiya4FJNR8onM2bZbahqPZP7SzhCp1Korhn34XLSM1yxBgAE
xPdNqFsXsZ2PW15t9HyitJuYSpuK83phEbC7BxPRBPRwl/JbA7Xe8CmET4Q1xpTQF+RW2M/3qN3e
FRy3zPkOdLc66SioLIELxwQItkdwLGOFHjEfIQE047N8fI18GyPdxqDR4xl9CsN1UynQ/RCc0x2A
Lp93ok4VFBrUs9d0zPgVCBXHioUDNSeQ3DCReb5s//x0Vp9gxcHqDMVXfvGLnLJwh3F8WUbVdn7V
5u6yLZG0jN8IKeb5bwTtb9Z9xdGM4HOpTxHWQQcDufsPR4KG2FGO5rS+SNuwMyvPi3u6E6Nt8GS5
9XBfKBSsOtpGIfWlo+FwZuLuWqVsX1qOqYEv/zACW13tcyV2gRCjYK5g3ZlUeDMc0xydL9G6y5MR
av898Wr6acwRVCw8ubNHCkCTssOKR/BmZfQX9mM7I0sDJUoqNQeyhh4JmeK+/G4Xh9d1Kajj+Rz8
6ZrymGPk6THsJANXEnAB0GRIh/zBe+yzj90/XeETO8TvCKdbIa2GMWphsUwbIpoP32dPSid8Pwv9
lLzkchAVaB00d4VFtp7T0VFZ8HCObUbKkQpOAZljF8hn/SLcf1vYj29wLta8j38iMugT6yLjpX9p
MXjMmbk4XXSqrxz5Kk9BY7HyXHNGGd8hJokD5qWAuf9oqUaXpDX7pK4hrcWw0XLSE48aWd4sCJHE
mEj5l0ZHmIbNLJ7q/R9EX4sg/0LYG0AgHKoHF+Yc6goXdK4IhJkTmI2FlTyl/moX0lNG5U7Vkitu
kVZP6on6GYVn4z8m+Zms0qXp8ckIr9Z6g1zvzZLQx83EE6ytR/UVtDr+EzUkG/k0GBHC5e7qZTtc
CugAiXoDLB6T327DbL5ASbOoq4pvcVM7nhvEj/6S2jrvSHwmdUwizeBkUzaoGXAEa3UYMV5P9yse
mXc7tf2CCWWnd8hKNNEph2GhpnqoaNudqd8+AOOx+dblUZ1lTIO0Dacv790tOQm2qIK/bxtO+vC2
CCmnPLKLYv0X77AEKAQTABsyv2wsSIqtdR5A3h7u7G0ieUKSbVIeWjHc4hl6YpMRpCwqDVZdQ+PG
tTvmMifbRWlgnSB5MmRsbBOzC155F9t+uS8B7iZ2o1AiS73NtRaz0r4ITbontnDznmwTbpCkCLJr
X8gzS65n8CF0o3iLVhj1Jo6adKAr6ZS/V9nWy5K5yqL8FaXVl5KNmp9X19Qx358+V2RVJj8ptw2L
K+GLVE9WhU3TSNHwhv8louydqO3UT5OiazIX6K7K/sZ/hLZZ0EgAG4EgazYSrRHmeO1gSU9MAGuu
vj/6fWSEIIir0KIG9X4EAfE+9Sc6bJSB/uvDMuJsfgGyL08O9UvpqVKYbxfltzBZl8WHp86yFqH4
Hhx19p+/eFLUmLuw849KCe807Xd/ivyYXRQ1iZZWWOwWa628w7eVusEc0kcltJLSGdzjPYEMDNeZ
LUrgcb6yS/1NIeerJpezBQ11ccrNs8xQv+QOExuw1G5qjr7v/hXhiJsZ4pWw7DtfPIJ+WooZbrJ6
0HqAM26TKdCRpFgehIu/pqMfltfSWY93o5cxxqCX8INGoVNfDpMkP4Dv1ZTT8PyDkd2m5ipTabXk
4D+QsZjTxKR1MN0TutkBQ1j26lYm6s06nAwqfkU3gXsefOccXcCxUVakJ9cgs/+k9+ccSL3Rtx6c
HVqKDyzrpdUwk9Y3rJYgUVk9LsNVTUyk3giGN8nnXzMEJD0D8SBuXi5IgHL0As1PwjsSYmnHA2jo
NQVvR8FRzZFHoaOgMhDtFZ5GwlzY/ggfagt9uoSTwBEd9W6AGixGV8W5N34f6CNmyQszlAMBxJw6
5oAP2FkZXLOLua4b9GEHZQu/mlgEnYFjAFgTKivyOeIwK4+nbrwvQiT7mHMSjhCGipmuel5uGizP
W1LSuiAHtW192YUFsC7YepU5SUkWv3pZRzv/ExeySdZfKpjE8mO4b1ej9ML9rS83ur4Ln5D4Xobt
dn/u0PQ3JfYP9Niqk5S0EYW1VIPao+EhRpJ9HjM0H3kMWhefYbqfDGq7+LyvU/c2zpudp7fl7yB0
f4al5qAPLNsXCxBNCFxd8SBWiY5SANleb9gRAFLRmYCmxpIi3Ol1Wv0SK0Hg+8uxsYKN1PwQ8aGW
lUg3IgXx7jqTmF18tzzX5MPT7ESOEEk1iyDqrQMNWQt7QwOtwqb9qlt6KxDwzsb/hY1qCkduzJeE
7MmYrGBa7KXm9cOdJd5sNWAw1WgaWIxvzEpB0XX5dHt0ol6ZbiOoMvXHEX1KNLljVj6AiyzvZ+Yd
OzkzTP661BdtiLnbNOisqZGLFKef/LjUNEDtgi9verN43wwDCIS7Slnm72M+nNr5vJe2mRXNwuae
dy9QbVDx+mkZ4yJUAqx/MVok3pf0tUhsmKMnDH9eGLOWOUpVQtiY7GvfnuGNfGDW1k9Ms36sx2PA
56YxLkXiDaRzBoE03TeuFfgTOOJcpujL15rTZQH0+EUYJdnsVZMW5Ty+fbZq377yKRypEO1Wr189
2J17L76p++Cg4uc8JmR3QlUixwXJOoj/w7uZ6swRoWZ4htzPn0onOmeMQ1/lj2UYfuy7ZjkTEq4Z
z/suj+S+wKx1UdVYNUsGeNBpIcF6c8IXpDx2YnOzuQcgSXlLrAt07TEvgG7hs4v6myHr9cVNTu6D
x4uzYg/oCUy0rUxtbKuXfRP+2ImTJSG3/jYdZJJVNiA6tnEFPmIx3eLadAFe4JWvar2UQsRNOPgF
4TqfYKDnXObPmIMdx4NUpIf8zLdJs1BXYmyBhdB55aLLp9WR+w7s708sm3/Q2NEJxg690TsMp7QM
nzG8YM8ChpoCL1RLU5466BdoA3rcEG/BFcPAcJDKu4ihWh5LZFWoGL50Mv6dDQU9avpXmwMv6aIP
+YxfZrFcXf84BhMLn82GTbTmBqcQWXOydJa2s5wzanA5AbRWakmpc0baBkrOtqOXan8B13OHsqXx
0+WVuup3uYzBeWD+XgWXQ0RJiOfULuF70QE4LjVfqWknDpJWVqz3OrLvwI7K0l7o4ycgU0LUImvJ
jeaXNg89YjKEJi0wAizvKAlUCZUtLALCpuwwpA33gz9NFYdMkPdBn+Jn7LZyAa4/lat+DInpFHDB
KXllKXqfFN2cZNcQ4paxEdcXIzQ0s1PcqY//rIdPPNPpik4Ob1E0cnqHIfRujYaisr96fJvDFezw
mUr2kleUZyKOoGn3Yc7PZU1Hdggn2VeqlqUb3Ep3X69NaZ4YcA7q9ZZq7oaUAH+ZChKUgl/WGCMM
+nJS951hA0P/U1Wfm9GJTmtLOu5kRIidZ0IX1FitRVojp+2JSUeUx2gvhQzx0bAV8S0qUiftCGe0
asyaVi3/CNmZy4w6zNKfUg2c/PAFI1QZXIezZdtkv6BuBNoVOsJBARyRNn9aT84MorIrNEdjSIq0
MXg6mkuO+/bvCtXfgeuYgy/pgLuFbfmQkazKKqJ+esXLne9sPvOfKvZ8pwlaFG/sZcQjo7zed/X+
MeLMt2a/CjwrZp2sYB32SKr+TgB6aFMbgBPHzBfEXJw1697Cl3QlBLwE9iZU91+6F4dCcLercYZZ
2WlE0gaLBf/TvNQO8uRQIZsaTHaR9b53DD4vBllsDPsEBgFT5KEdxVUU0re4UUlKBHOd8mKX3ZpK
VS66muOh1FNgwn/6PyXZWQDUdSN+C/h366DrFgWLRWvqZJ7sKqLCgfGZz0VzwjgfBTwJkQ0l6GVx
H9DCL7RdbSbBuW1T+K6gorm20IPlhS7Fkl5y5jWMFzDAbK2yw2akIZJQ73FGnnWHnEv2UqYoatbI
0KZslrDy+JfEXkqR4w3S5hMBVaIt+3BbWYtQbw3TATpR/2EY5OMHTtP5caZ0Ed2OHw2AQ6sA9zVc
6EBr6NGKspet5Cg/mWs2I1cU5diJWzxo7XfMrIA47MW3zwkce3cDqulg08wVwqVoiBxo7SeO3JuB
MwS0XPPogdDYBz2WUefsPP1SN9/QjoOWEcNRUrYFmYxHiOnrjBzx51Ge/V759NYjCWNflTipJx3+
JzQf01DjJoBOmh85LbHnptDjotq9+2S4J8ELkhxxWK/ZZriIO9CkJqGfofRSUtA4yfH8AmVJe9HQ
NpnWuwl27ZQHX1pdTBa6ZN0BdMR5toWd+40MDjI1KVfKZc5FoNK+hQs3PBLUV4SErvMSPKPigei1
gPYy64sI5lTNx/jxaOnyyEtqKNWnQzP//0ryP6S7gqSMNjYMNJsw5bru9sdeSHSkPLbEeHXOefpz
vv8v0XJASAYcSjBdOLQCMxFJiehqWJLZ3sAsPeAjUwi+SQxSlyF+iGXTsqRo24A5/LNJkRXngH7N
lbwlDuDnkVU8oA++f9BbsoA8SLLbu3W6tXfTMw+Q4WQp5f+uwvoLWtOce3FSyn8+RsPoL3D32GB8
EgHctRFZH/5KeAAd4Hu/waHc5EWTiGZJMApJ2Zdir27xJ668Gb6S1qN4pdBltNuUJJ1d8Smp8ZdC
aXpbKX8vzoTG1pSztJ/NVV41gMQlDhTdMX1nnn7uLEzJPuxLmSYjvDzi+r4OQfgQ2kJ09GHXuD6B
HxDrAXSZXtvnVGdJ41oSjWEv949iIUODk04qAxaZixRass9jFYmx6ftBkPLVPRkns7ayvk90vFtk
UrElJEdn7fw+N40AlfW8M9AkfmnQkKtg2OKGwMj9iahUeG8VFB+gHtDJ+uwO++SotA9VWdd+uKWl
M14pFShw00mjC0b3gZSBQUBjF7tQH36XxbLzNLM8mHF24DB69TU8KpAUCbn2o1aQfIRSISFI3K3/
vaeogwxLrqD2AkCTumU5eTpQpSJIIggYahEE7ZGIIoMSJLVL5YL/+nBeL5G3LvbvNbADqHsqLC+9
VfW5v8uOATVbV//BeRcnEL9D/CcMVkwjPTjqSCBG8pEKH0JyiB+OEzr27YgrSXJetqbCZB4/iCjA
kbjH0fk8Eo1W8/2M9eJ32HrIqQs+sC6DK4b3LpGi+KgQJvPxfEOqjBeVeX8M5PVphZ8NtjEvMPY/
jZESthav+CVOo9rroXWfJYQ7kz71cu6Qlz1T8H4j8Xefz3WIaaXWNJRmbolfk5wPM4/Tiq+KWxIz
2q1s/ArDK3lV18GLWnH0CYEwdnRGkEuTI6U0Y95pCodwsAJoONaz/BHl/TYOHfpd+fGCxWya9JrH
SqflKlBziqmRCm1uGbGJPJmZqJDQpX8F/6Ph1nlc5s1wp67LN30bOVvrO0T2xTqmE20Ayw2+i2R1
eJj4RpcYopNnCBosVMOe/sMPwGMkPy0th9gv1mZBvmqvVgl0/Oi7f6QqSVoixtSPGkijByBd3G8u
JR3DNTymj65UBQKWtc599fA2WV/KxtCD0sFA7xt7LQoMFMqbZa7d1ebRmkh4nih9rSOp6uYJmFkz
4NquZc2u2BcsQAy1m/FHzVZP3JARPetUGYJPIkf/BzY1UjKcWw23JcqiEIi8llKIBSo21Z+Dvu3n
BQrq/tJ1sbOil0+ibmYMWwJ4g3NKPoTTRxOXCorhQqwRJcq2/lNEisMmS/PaCbaZNMOYKmBk/JPI
thfDf4cz9cEIF0in9T1E9unHS/EXoZ7TshZb6SEDjBN19u8MkiYK7bULYihPJfIQn7mqQcQjBieO
KsAmufI6get10GSNKLVdG2k8jTFDCeQhS9MYb8D2gJ7Wicxnd5NvyS6loQ+rRldxuQviBIypMR8w
nm3chPW+rdbwBZssncJrkgb0U+l8/ipXXkbdNDHzs0vxDwG8DmRAZpuOLsD0EjhLDPsBq/zzxPBV
u5KFcXdLvpgDcwL5QIOzYiptkUxD3CPMfCMqtS5/vagavh36nE8MfDRZA/Fm+PUZayY+Zkq9E2Ov
mF/YaJod+u5kXRL7CyN70sJ43BaIto2WbgRYJO6UgoAiNR9VzRLfnJ+m+bMTQW5xBrGBeeCpc1Ba
xsV5TZXaJJKCGrPuHWaZFOQ3x2mlDdz11oD4HHnoOCkkp+WVv214xr7QzEdRc9qpal9kJ8PoDLTk
Iu8vvUX5DZqoyMHeA922lj/k4yLjKhs8g5lgnzu/ntRuXsiI2qN7XAiccMDvmWVxKpnCpElJaOei
t1fhXnnx9UHflbN8Pqd+G0h2GjC6m6hpZMUmWWkfYUCkXPtesjMxzokACZ6QHHy+vRBQrqHYbalL
nwe8M3ncrRsO/7MOBkHTRZ+DMRoParDRn2bt4Vve+JUVzlWirQpyS/emvN2QtypK0ZN3BzdjJ1Cz
32fIiASWX8wvx9XDn8K5xgzv8HzSJrbZnDGz7/KBIY98Jw+05+Z1eNokZTz/eCDm49GY96ozSyRG
hgPPnXvHkJ0yEtsP+ooO3ry3rNo10JczkniXDAsRgiwv9J/zE2lJedHHO20V1qeAX7ayr/Re1neR
Km0K1257yCmxqYL3KZA1f3Xr8o+zYCaHGjzjesUACdzX3BTDAKlGtflfDnYOFSARGrCVpOObARi5
K/b8lUIP6DAJbMyUvdOXH55xH6yQXO1p5vDjVo4CM/UhRdwwwS+xCIg7dOw0RCeNvx3OQAaH46HW
swXcglS0wrz5QVukkZ4Tbnm/eu3uFxRBOfdvK2HF4+uWZgfC50XOynhr3N3Dp2NmH/80I6pyaYi3
HWrLTzG9O743369nt4Ak7chG1hnZNHXbsZ3UX4Pa7o4wL2HHZ29fuHcsD1s7vZNxFduBkMwpvd9X
xW6aGq+XY6S3BtV2rxmue0H9g+xfdZJYxOXj8O0uhJKR3s+GGmySXKg4Zq1msaRiOo5KJRUIrk8q
M62G94XoJ7iS+8VmBsp9u3L104N6lb4ESc27KfMbtzcBtoieo2F/eAEcWWvJ1pUcZFKNsLRNI/PW
5h6cZBOcRNZDYa/HkijGLBA0HZZ03ccmeHMmpPJE5sLTxaemCLMc03Xlnj4xy9EBlVj673UIgQxv
HyLuZ1Gr5fEFN6sDgUViL2mCUgcsluFTN9Mdxqu6DF9+tMX5Qa2t9LlLp6TGYv6mtjqlH0RFsTrS
mLOVnMO4QZx/UIyuHuhG+M7pl4guhpf/F6XbOIitVE/QyHVm0aqDkhzFY+/hGDzkaJkmAgl2Pe2t
W4yg+ysSzoddDJbJeopCRDMC0fNEJsv5iBm5lIlSnd+CorHQT/LZCK5vzcMmuexEJBLj0eul1DYG
2x7zRGA+fePmPtlmSRQ6i7AiePTxkeJpVx32lGE4oNk2Ixhnow8aDTMQJPvay6KnIbCZS3olCWWb
zCCRyasrRhxHyJ7Ir906l4ZODPFHf1Qhse0jjYTsJFC6vxSXVpagK2rLsJFRO7N5cTV/UpNYKlUi
FoaT+w8gJKh2e/IVbR44OiELd5ipoi5c4FDp1IyEGbqZairzTgrEdJh4MckpCeKNaIw5RFNumLOh
LkkjzFxagyb+sKxNTmIzqSrE0pScwNnA3QxfiEfFwUNlhxUWPerI9cqvODR9CtHfMPBgdCigJ+y7
UTfS74vUmzUASwEZtnmucgd6YbbjpnSHw9jqcpcR1uddEldZkayUeu0geIy90e3J8T1s5KDPpmVi
U4RncPf0P5MX2Wlj+tamEOCxaI9Cl8O2mWbNaciSt1SOIz7lN+GMoVSlkCRpzMAdWnuO7Lypfv2z
TxlmSIRk3GDEPZ2xjaHbLniCr7BvlYEzmcYlIzQ3N24kcTsjKuG2OU2+jUTXuZsrbdApft9oaPP2
CcJ1JfJ/OKSqi3QjVnCdQkXXCU2N4/Pujra83ienlKRFr3ymWAI8H4nIX4zm6SuI/b3/ImCh3Dm6
21RMODGBvm4aZiJhW277xsutavrwz1BH6xivcdnxt9q5+eOoG0wIIbaRy3xwsO6UZELKLSAWsYB7
tja3N3hRcRVxV26gIqk7aQ65TuhKIelRznaIF91dsjKDGJRnz+2TSlwkTLrXCabnSRcH6k5y+61l
um05FVy7z/c9YT+2t87w0JhH7hSAGh4wAD3Vt5O9oOSJ0ZL9OfZnPvt1dBukOzT6JvmDU3LHXzJA
zaS2Ge5f19R50N9VPB9ejXgyFU3KlI6kdg/eTs/xfcspAX2Cfq4SzEgEB7BFBrdzNo3htbCb8Xig
xKxUD3dFO+ALDY44IFlXGFYcfA4GOfPkH1YfJ1pfBGsjJG2eNeO/y+vaymolyE5G0sW/n5foS7kN
lYPNSEjTeq9E1A2WWZtdKQx45U140MDEqDar3MW/9ELRSE7HS9j0+dvUwk+O408B1i0Vi1s4QsdQ
x5ADLrenu0lK3IQzBOqgFqufntW4nvf8M9feuLjVqBKIVMOBLW1O7c30Olq7vtglEL1psy3CSDQc
CejxCXwpO9fKgrncXUM/bGjUe3wjlVYvMxPolSDip5YciypVlyM1lmhFRgFTIkBdk7mSQpOu71CU
EdmgpYoluUhNjGnemp88OQnUpGC+i9/IQkcZBFso14BXiEfuU5cUxwLQ82CsiRhu5C4VSMkRLlv2
1YzqBMoI9MVgaZr9g0MtK0FKh4XZKaNN9n4RQY749iHzpqciSjgbHlqFKii7J2SiCc7voyXXIFve
Bo7ChaOtSomm+dWd9hcp/eXYekqfvh60z9UikU1LPJtVXkgZQatj220v6at5IX3bqLeyNJBBvcg/
cDHyHe+GHp8Iy47XRbnF1+xwb5YGlX/ZEuuLYo0rc0PrJKQadd2s1acaG5L5b7rmSKSsT1UUr7sO
xXIcsMr/Yo+MuD3DiKZIkZ8b5Fi2YsrOg1zeGOQYLuimMbrqKnTeFrRaTHGq0KitNx8h7NNXm1rN
JS+Gp8qEf1Es05PE37GKVlONC/QTHlDeh80T3BBAAdNWXQRSc04+7qHdIqbbOTv4Tjg8jqSnyA7A
beO3y/k5YDA2E9ZHjMjvo0vAnKbIlVv1/97uM9SQhtC8jRuqF6W7b13uV9KgRd5Ouf27fjroF334
MOpCKRlbYnXGpGTos8Omt0WFqDgjoinGdAtOCUF40VquQJkz4yVgGIrA3A4aDnSh7RcAJtb6gQt+
dubzE9JTRGziPskd2I+FYYF0uFPqQ6P9uyL2NKNZGonNrzzny3TBGe90furNJV9GQO+4uGmokwAF
6nbyUbdGK3sLuOrualntKvvoJaXc35JE8oEGZCCvuE3dQdjz8zq3ZI27GNYmB3L2tamIc/MffjhA
Hka6I7XvOJkjhXv4ckMVVXaUy73+Tk/tBs+5UqPazOv1zFLxDwyfsGyTjMk0f3NWks+STwYpK5aa
8G4P43uY1GqcY4RcS2WX3swu2BzYGwLyixUFHzndxMWJ9LScZAYB/L4W3+BraZcwkLJ1jZcUskyZ
dfo0juP1dfirT+ofbMJds+q3ACdcb3tF2doUiLlzEvDUseuqhB4nbsO50MEYKNn2LzsTHzKoNTc6
K1UJfBpBYilZQsXjew65yMkcWf8YR/uf71apHVVmtmwdM3AtJ2u4KA5uFg+edEaHmMPa3IntEPCU
yOpIiNLzHc7BcGKm0bx5lc6wjIVTcQlplTMddrK/XHeH4Oj/8UKGiKV9LOAxGpRY1viTF+NGKXpo
7zSnoObOx6ZsArLSXoi951kpEebLXR1ZutjqTC6Sdth0b3/5mY7PEmBNQU5F8WM9I8L3dJX0M67t
LOi+5IrH86GlZCmrJ3/J6SukS8Hh/sS/8GZ3nP1SpCu25ZpvML8F/HNBeCgl/ZkwB+AdfMn/5sY8
FmlcjGfq1xPvfce2Yer9lOw0FAkeIMuQYQa3cvpDTf2tp3r6YOJ7nxNYNbCJSdCz0Uj8dt0LQssh
v8R2a94DWAnRDqORbml8rDTMLrwFAfcr/CKGKf0c79Ior+XgkQdjXN1LerW+RQDfZqBMMlj1PVIY
t2BCMtfePapj9/RLRUgTTg/t7AlI+5V/hoj/I/pdcek+IEolXB0PrFSDSnIJLjpFzrSX9QkbtICM
0vwzvGm3TyBctwbgGoGVYPMBy8YfdPJWfxf8wNVfBODnEEfct+5UUmRost4fM4TzZIPMGRIxSk9O
2FKsV3jin08C+XRi38lT99+ca4lsgV1ns1yQ0Wc2+ttsYbXEC1/a9fskIbBqrp+xP2rW+UwmHX7J
yEOOAJR69wls05wQpOqmmAUngu+5IyBAFIjkPVHkf7IszEaisaC1/mnlt1nGBJyDS/GGiXWNEicr
5mzgyieFWZuIAAeajJa+6FSkeImoVPiWuM1P+PoCXvzFmu8oeFdNW1e0vo6FvwfhzB+bLSKslMQ4
DIDn/AWs7hXgABM4A9m8r/ib7ylgyrVxLIhBlod2Rjnq52QtA2nL3ZN6wRsUKtXrBySMDqRrfgk6
rKMPGC+5FNq0bkbfrPxZb7RUV3oaoqVAE4jxs9AzOFWb09pc4eg5p75fYQ2y1yWt7mWYz8SgIZpV
u0Am5b4RjqRU9y3KGPwkJw0oNk0johO7CT7xOF7homdDDCnOQUZvWzLD6ktLHgmmdU9zQ73AvlxI
vPYfa7f8iJZgtdGdWGAhpkRXBNtfcJyH+pO8ZDdNFPhEeQWqFo9uGJlBQufxc3EdkFhp7GGiFszU
1qKYn731YAcL7fRWbWgU/LMvhobCTQFNYjWZVhI0rm3QJDKaDa2xb8u7iLuPwIOYQI/Ek6Gb+GCQ
ozbNaKP7OLFFx576zl7rZSv9EDcWDBgqmJICy+km3nOYLUgVytrow3sd6R1yu4BO6Cw2lLsZUXrR
A8KG8swtFk+AFhPxDqsi7p+Unb6rU/B8qYRFhUtv0um24EB1HdEeiyN9KnIKOc6+4pBonBNze6eD
8rVhZhrolusnEksbvgd5+2y+qlyFN8jsIwVydHq/4om0g2ka866X1TugwZjFn99qhrlP4FZz2R7y
QwajcY79I/ehb9ZuX9suIcP9g9mV1VCpC07aXzpKv8YjYpP8/IuDIOSGTnanauR3kfEQF0N/l7Ig
vADrLEE3BGhvklmE7ChOxT4IezQf7TFPTb5s74x5kqa2sjWA/y7/WvlAdehHqAez0v7S/Tu3ZcCe
KmiXYeUhM4ZlEl00gnBSQJMXPYu5/PeR8CfONsZsWSKRVguTtED/ETLxHDZVSgr5IYnIdPn4Sq9E
0b/He4R7t37pRabLul3kRwTKebrQEVmgtGv7xDnGuX1l8AFi1T18HOLdHiCiJDXrzMce3T83dRnW
vPjF0cyPmLJYhq+0vmFLyppL4qY4blwYkDJOAFcCdUv5DomEruQH9qqFrWTk38sbunC95y5KED4p
LdLTGmth3G9SmtLX2I2HO5FY8MU4ADccH0oTwhWumtc76CipbYaLHIwGUkwW0Z9nTqSRgVv9e8+u
cZ14j7BH2aNhIFMTuRVnf2GeMPSXY2btXePslppYUsu6jrLAfqN+UjmniVjI2xAj7sBrC7UflldA
IQJSLsQh5jV1Q5lzhNlK07RZJzAGoIVVe6sAMBil78SAxeJCtoKtwm3a0edXJbWclSV2cUF3pWa7
82zm3pbnxnPE/VXPirwV9oG6Pw7xfMcy0k8ECkMPx7apmrX9081FKPQSM8L3OPixjDntu3/qzkHg
tWXI/kbvBIm++Z7DBtfmccPlx2E0zta8aPgF0PMlNOFQcviLeyBhVh4s6jS72hORaUw/KQN6Bx3U
6Kx1N2i6M1IPI9UdJ6WKayXKFL3pYUB2tVCn3yLduv/EluHk1f439T+Ss2IGni2MkjGWXgCpIO99
FYyTWNsWDu5j8y6qhCKY1Gp4500tN5zCWURzNAHs0IFHBdsZ4CHPXr0BvgGxiS8EP/0CTmjOfuZT
gNypk8tmXf6bmNIxDWlGxfbE6AWHLQUxBn7X3nTMQLziOpf8oDJq9uWEtGVpss5RVxSoqwWON5SF
1tchLENhTPuP5q/rA955hIXKdXzbE6/M/U6yr2tMJNkjtuoF1PzZo6e+V7DVOPCIpU09/iUoB/lp
ASgeHd5bL4BU1xpPBkG5u0jzz3wO8wovTG24/nKkXLIKkQ3jbGfB/Fz2jswzR/URGc+HgMEVEJ5m
vRvgAbXlFWlAiHFNeEuyu741ODnPR/pP0LgcUdFA+nyOScW/nLLu3Hl/a6K1cbR96KPVwG7XYhtg
20Rn5N+5m+LFX6eB/nxUSDuLl2fK9pNSUPCj6+oMe7TU6WnU/oJQLbF9KLIFhCRmsp39nYuytxaK
1MCJ6aiZRw0zEclEHdLxgweMkQpmzLRkKHrZNIbDB3xhIdHz+ZdkPGbxNSgqkK3NvkxrXZg2GkKp
l08e+WlTqT68WK5MkgXJZyJYQwGfgon62r8BKAM32kArhcnZX3tgZioDfL1MBpCzoxZ4kLsGVHD2
FUm+eT5N5OeHsh0Xp+fGO1Q7+KxB7+IZ2vjq7ywHmgtHtPyIcuO7Izfi/LgEoSwAGzHkZS1CZiUP
sOuntdbnN706PVTN6UifmvZu5+o9/dw59wky8DRw/B8/tsSM3QI9wKzUWk38LOnzI0KAiI8wrD0F
ydmv5nWju7HJ19kVAyCzrRyKh5BNEVbda0xJ1cp+KfY3hqVmWvJOGaCiNMrDcGmyQMcX2IEIbLxB
pTje/rc585/854QN7gO9+OHCMoZ7kxWE+MKJZnHiddn1udBPTCEBBUMRdU8FFyDTVGCoh7cwsqLs
HOZzsQNO+zQOmHegyXftYSVBVXEA9cBgAKV0XB9Dwd/8lmQ5SDQHpb4LrxRA9sDywhH6RgZrh2eV
0QVPG9JvyLq742qxrhHQ5CjNF1pzd/69kSd6BjvYStrrNFZ5WMoJ0HWVUJIppfrhPB6fO438eE47
dqow7FcNX/a2dD+O0kjOBYJULxifqzpvJreepFJIPSTYUJ8D8ucr5qPhEYBn0kO60f1HwcGh2mI4
PB6mVodrqwNoxffbZnKuH+5GBrVV09mI0xfMXSKdNIVN5iEgS7MKItZftOc/QYObv3fn6puHW6Rs
t8f4x+CyugdxL/6rSfCUgBt2YJ2d1m1POOJuvsl3eq/TjpTSftGHLop8K5q2p+PMTWjpOWcNpi+B
TGclIkud69jUh/TCKjRumrH/WhDIFxpLlYfx4TGOI7+UUtkSqiscJ2pkBzLxe5U2mwvld9ckZ1eJ
bRl6vtQQCSyb0uFZD/GN3O0v/stWJR426lSBJgjURmKDA4VkpIYATWqvOeGVza0BN8PCIrBu3mIW
/6UGtNVUPq4aCeXrMmFEkzMLMtajKDv3I0etjoHXyTaCw7a2KnA0mEleJHLCUZWMCkrDlG9eJQ1H
8eF9eXQZuio5C/ArCUvDNfs2JLuKvQjQqq7QfzM3SFkGEJ2YG63TbhUTXnsHNK1erbb518meGvyg
cr7gPqm2zgfWKrBQ8cSU/z0VNClOqHQ7v4BE5AuF+tNR24TX24D4nHQm0DuMqX6WuJauXK5L3hdX
91kFkb9x+FKQLZThcS+On00KIGPRSNB5doIDhDBJuA2PCXCKxWMVDutcyQYKmeNVdzApx2nJnOU9
w3//2d5yC8T9UPDqAQUeteL5UT2jvUGCBjNhW2DWN22ass3SFjhLCA6UkIsdzg0QS8CJJUWkJvj1
wd8B7Esv4nX25tL8Rd0p41ft0ChrhXru+CMOxa76inRjSsrAEU45RjtuFCPDKZVAear+3O76nzCZ
1CiU2GGeZWzjodIY1NQw/zCVPUrWLE3ZDL+u2jXO1LyC6COVEozuXE0QJndydCk+ppq88PJ9FFFX
ov9WxwHkEnMMllTp3NFNFCtwsTNVsTW/xnrpj3bpx23cEX0Bz44fq0oQnQG6MlPd7dfyUKMZElti
Hg+hJHz+Xy39fS6eWKP82Ng+NxF6UQ9jDBACNcCAJlMQEouZOoQ3mynGiktMhM46UmmuxX2DxOX+
3kHs8wpXFfkZbYOJz332s4M6FNGsXUMx7yf3dW7Kxnoj3Wm5dZZpZUDQfYRY2mZNu7nFyD35qxde
Bk0wZAeSF0ikkV1we+0eZVpTvmBaZuIhTBuy/UUueiIudDQ1fWWZp15+jamcYljCro++wddg5hnK
xCqXGBmJKVJVGuPGMR+tb9VbAzM2eNYtiWEoOUoMYBghLRB46UaMU8n3HCHGqLzbc16Y2idwtfjj
3YQ5tONJx7brdYnXxJlq75vLN9/0Er4Ry1X6j+AvqYwArjJ6Ob/L2nHAzQbrmopVxJ31w32dTO8y
42/eqIpEgb4raXZ+N4fHWxp8JSxmm7YP3USigG9MJquMz72WQiSLdBwgF9boKYFSW2YNp0feeyqa
13eHiq4zWYsyTMsQymRQpEA2aWCWrV0RwPqD0JLFqBcp1iTYjQENehroH9QjcPSDjhfHseFrHfou
ro1hCHQIAqyMfdmFaX6KsqAjNRj7hOKdwxXa5OAUgrLMlkPCDuAsSWjOR4KqYN8nr4Ctp2wtx80m
rfUlE0VqlfFw8+0gayGUIOdtvnk5kxh2hz3GuGyMeEP98ghHBlbcIzM6pPo0uEjX5lE9zGdvKwfK
qt03dVwNUvaMD1IaZioR6pw8iAibcS+cgWGyG40jR98dkHgtxfRga4SleLgjJk5KabtybVO4YW5T
NOh2xA/WOPExfBPEeCQ2yIqFzJbCPFNz26D/rElT78z1zb2ixm7O412Kygnok67mJAOHclk59hHR
UiGX1Dy6XwPmhs+ie5w3ny5LrPy9UTVa1UXbYkHa3A6GH3MDW2XRPBXG56hzEXSGPrWqjnhKyQSr
/rd80f7QfwGq0jyo5SQkVTiqXDnOBjPyorfo03fbrihfv+a4hUfRYBM9vAXhtXJJ2XwgeKjvKGr7
XY9sEENDbShTn+isPgcJ/OgMeh6wY0Gr/aYy4GP9ts6fgkdAzEamszzIgXPdSwMHfbj8er1WC+Ms
HuZjjbpLIlyINbHhU++Mb1FNKAZNwYj1YXUd5zrmRBZVnngy9T6msInuTejh33pGsau1rU/0o5if
bmhTk67nIgY3X9LO/TwWWNQs0Ws5WANY0xM8APVCZCgmQQTT4HRk+iV5IDcy3R/+neFS4P/xtrt4
/SNd5Sm8D2DbW1LJv2Tl3bbcvjJKUhWzFDC6Dx8pLSKgA7n2mXvCwyXZaCKtba2SygOk2AA6+oQj
J3LSYJSIKk5SJ7INtMhfqzZiJcNJkqeM6/rDU10wnkP5XB2DbT+S2OoomBuMJ2lIT9NS+z0UclhR
i7bktAukqWPAKrizxwNmnohKRAF0whYAEWIr9Y4CyMPMSfLgStpfBkPWHRjcYarD8UZS7yKVmgoz
2diPjp/bo10zelMdkrYEFzm7d9tdmGbHvgnAvxWZ9KPLLYmU+Nh+ZSwTy2YnwaRfTMnFPw87iz5U
1VurUxJhkFugEdKIah+W6VsZOo4PWBp0wE7ErDTjkxEkSEPUFKbSKdMzCzEX0cLtSAQoHKaySfuq
ytUbTiGhkDPfkBip4OMISn9XmZdRtu4tuD8fxckVzGFpewuGsUnfNZaNcy3u+NzM+PwgBccamxf9
3jKwwBCKUVc/mOYFMFp/RbJgvjO1tGRUCLvrhDNLTGWa33MA/Ej/Y7v7RBAPEWG8pGaJLWtht7kC
Abif11GS4Immc/6LYsfB9Imo8Jusk0xJk27+V1F33NOW5dFFyyZ3zQ0++gZdDikvUvYRMoEGe/14
uuX0uAhs2ykNnd/KWX2/AzBHgiSaEB8RTnmpzpnhJ8hFh0lchsxTRm8i5JwDmkgLa6lYg2GgDotK
3GlWv4EAa/W7Psx1Y4qDx2c+HnPkBw81gutadpg0yeXWAvCSkgl1vh3NvA0rO/6686PeaOpsiVSw
Lgamv766WyYCAyr8Aw43Din014zJR3jOmj4fkKjOSyQd4skr/EG+qqE3deIHrzkFm84VcXQ/d3S7
2rMsOXejfOtAQnWhCcEwcJDmW/Zhb1tmJWVuxueNTndqO71N2dWGxHn3zqw2VQrfXeV1FRNwHPgi
iEYbk7fJYPohAaoPrCz3N4vtfj323zOksOCumj47+p772SCXuMvYBWJ2VYsevmAdOqitw0tAxYka
u7TOxR57UWTvBkJhbjYITaVgN0UCor8gtPgMeJ8lHYTeRy9uL4e74LFnsivF5i0r60RQvhvWrR/w
hFlhMEyqfuwFiPwN4yfV/GSZ3BGGGYEBpWpaGIQWhM6fk3Egf5FGfhRCLtbIqNFAmvEK7k7TVCUb
DuF71kfPN062zSaLIA1u92mch4ElqPRasuFmlo/aE2+9J7FPJD8ezoumW+9/rHQQ9oCOHyh5XrTt
hN75tJMQKj1ZyfUvneS8c1AlFvcpOpPXrkXB/5pLIbi0s6uvHamlymwmiq9ras5kAPS0DR0ym/BI
ayLY66k1gYS1pRANy8g0mydJnD6FzOKNvKIlz4HoUTALz7mVo3WZleOI5MEDjRmymela4qp2f3mP
BHPvZ46rR56hrst0goju2PI8Ss8HJut0M8jV4UcKPUbp0NE/g2VZ+r2HEJLIIUeNRHn/x0Yh8vT1
ufg+T48686UabWtk7ihZFNZNgTgzGbUfWfE37DiqERq5iBd6mTGcoAGKn05GHXTBVbzH3B60SNdf
0LQidQrBNSPQOhIp3xy8q7Q1NJrnlr2I5JPrVYJnWWJOYNGdufZWznmd3qJkLsD61HLyMF8y/9fn
9vzBOx+0DVsXzkAFJlKgpbnd2PyF1fxPV197mXAWcBT3S3QERDM3bCvAQvLMjOJCoyhjABllSArI
pjRuQrhnnU3YmfyvTneCEQXXms+0CuYlSkPegivdwQGglmUJ1D0tsi282rJUGF5uKJo1OhVx4ofP
fdLu4bCDLVUQAMVDRdsueCnLp7dXi/bnj2pyRAeA9xL270B9e7ETKWJmPxLxA1q2MyH/mRfDOS+x
sRzzmNSXvsxGkJWO+1DmUP5rJUG2W+Coqx0W0s7t97p5HNr7Z9C50Y8ddhEQaUoSdPiYP3rAMHPw
MCYrXNVuFEDYwZDGhF2Rjrv5acKKkL61VPZ2frIIkhTapYapOzqoBydbOT9gt2QLHUiRh1RJ9V/p
ts+9JpW2vEjiqUiGLh4cfRhpKBQhQQgaBKOUKkPGOqqnt/M2BQEo+NuL4hUcvXj0YCc/0sQUb5ed
7Px8hEvUHhyx4fE2B6RtmyBI2T2je+rxcztcPppMrj869/T3PDO/jSYxRvrCxYaQ/taHo6K+bSiH
12TYZyRut7oBJYval2b1qF+AmdE7ft7G67PUhpGG/H61OcXUMKcIzPJJySgcj0ihpJsP5MN+rNVh
knbsxf+1LRGFCAv/D4KslGNwdQB5wdMrUDP/6WkEwLXMZibYUyYT3xzqQ+Yv28GapsmVRJKeyFpJ
R8qqWJ9O84qJ3LA20YOQxJZJsGdXWtsEin9CC0jsP8hdU94y1c7MZrqOy7UiALwD0MRtL/kax5nX
Sp5FPTmSCy2CXYM5CrGgzW0O+rw9DzdCM7hOVSYW5eWomBEi9BnEwXR4GPVL2eBEGSlqTO4VlimG
JqooMigVj3ZIJPwlhMX4Vdl0fQ6vQ6guplAyF/Ep9Ii0e+4+t7MxXbluKsxUu+0xEKx3ldHQNuIC
+Y2MtQydgjTLGKeBi3MlXlWU/m1wsUL/slsJYLDiGbEIVGW8tGwC7ywlSkwDtc3EqzCy5iONCFrl
YS5GiJ4WCR9hKzN8gtBlgVVPDQhNncMV1rivgxviB0RYaV7Pmsyapeb/zf7cDsjEaSsiA6vKjkzo
19CyPZgxYJaqgmU5QaOJlc92jYlonDP6zkvMCqo0xeNmGYXzcChhL4LcYwLCTrwzQMOruykVYUnq
zZYGfSrVhBabyLhNBGk89EJtbQQMJa0U/mxAAEM3IV15hZFCMw9zYW+ojJTINn1zGyd8Nmosf8ZP
lInpAer+mZ7BBBMeD/tqJKpIYEPVZ2XSDy30Ts7QT22xYN6+ct4TRCkA0XWx6tqjzw5xse+AGkVJ
TJ9Jry2M4vooZdLzrc7GBA4w1sGcezenSLN0lnAv/sZrxyyRbnXswqXjzADjFLiunT6PsVqCHrmO
rL0aW7Qdwct6wA1g35rOnlrSaAbpCm228HYn4IO88Jpbz3Lim1Fj8MOn2kI4VHGw9jJW/s1VLM0v
EY4DADD+VKdohUJj//rOZeeiwKjseyYyH/RJMhvQ3NG/oiFyfO1ORGe/IYqPDShdaxsHlSoLbhao
nZla5yxVmePVj0u2TmfYjArxm+rN5h2oF138Rz31aU68nLVRSr7gYbcrkcSxG6p7kVu7NzgMu5hB
CXJToUtM5JV1MdouDHDEeXno+Ek0H6FTHW9Y6tawRCxqr+sYj98TK33ym6AGO5Zf27Esf+lIIGCh
eL+XlNHDlwcq5LmcjO4E0O+js/buzQi57bf9jUAM5BudHhKXMlvbfxMhdLuT9Uhjz494d76JYfzL
qTvZaRzilcDtZ/dfXK6JBqfXtrpQYCqdTIcV/8/ZLW8QHm74ct3GPq7dK588RcoRLq/MVWC3mjQM
WdDSlAuY+8fiAJQuqF0fcNSoMx6TZwpgmqJpqJxBw0+gCW+Hw+Zdv0hSrbUEyqMRItZouAjta6kh
il/OmZ+YiguO0lKidWrgje/W7gaslSPty7lpD51WoDNIDK3R8pjpxCXJF2RJUE048+uCLvaeay0C
wA8pitIdzSoGrtpWK4tdgWFqy6qRoUu7hCZRSwhge8RqyDOlRAVZyyRtwoOLDeXe0Ok2ek/ClNbl
UeHZVRpPflj6xm3e4YIeC5gKnbRJD9lkvesF50BPlE0CtQHAP2HFG85MvdjmlRPhwgz9uXhAeuXC
j51ea+fIH4py7yanwe7rTk3ax5Nz14jM9/vsIxX6QUYm+lbPzP/MYcwUQG9gt93WK8w+0uSGS2VK
vIVOaXyAewMOz5IUdo0GbuxebRACWvw9A2ADXDflbGDJYhfWjoT5d4lUgCx0PBdPBEk9fnerHLGG
FdiDAdwP38By354qf3SCZh9zDqk6hkBYxv8DwBf7IErR8pmPMc+jedWgnc77n9UxpF7RV1vzyoCP
YevW2ROjcBqw/WG+J2AGulYW7Eh9Lsj62Hi+C6HaZvubgNHFdalCfd50r6mTIPvanULfikm2FAtB
ROj8ID++Arv346L6hC6d02f1ujvBhzV9f6trPbz13B43So2p8EKqd8P13JI599BOYT34v2R09HfK
vXNIAKgEykqxWfcsxRpcePqT9PWAbyeR/mGsvjk5I48AOvU3kVucArjC4C9EDE4RRH3JQiFvY3QI
cxeXs5t/4Z6Xrg1tXkWS4mIafOTVpqS5atB2cO2yiy4RQLk5K1Hiy+yUVkiuBa74fFbOTGzA1xc1
42tt43pnykmCiPv/BqHRCaRMaz4bhwGh1QmkEq1Wiyq5MiFxUpg/rSedr2X5Y7R04Rr0KHnUjFX2
jsajWHiVPwkuXrtOYCELuuFtiKv7Fc8QxJpkhY5OnmXYoFCNTsiL803nhPHUE0M/EXUIo3vrsRTb
tPKFuGIlVAnNhjKKvY9rgIqcSvm0xUd/I7anJaZSVdcjO9kLvn4Z/SPdCRsNN6MwDoPdkM0q1Ehy
6IgMrgWZLtQ1kGxZzQTI4nXjaZ9j4VooRn/Mx5nz6JkCfdzy/sk7ZWvGapgQ1Z8091sHqfxl7Vkh
4mGKhuOVMK+qCWNu5rhojdC6SCFBUy7ZrRObiXlozrjyy/Gm6r3rDE8rnNWYPHg6WD1hK+W9+aO/
Esbq7WVVq1FRUCZsqcv4QswZT9cik8cD7jtKIWpbjziUMrIh/xzXfqbOcXFxBuwBLyAkT4PYctxg
RvFAUPJH91aO1b6QW3/t6ZCSv8bfwqyRALJTwFdGflByRhx6r/dMi4bXiuHl5fHFkelblrbXbwmr
QOoHPpJXtGtrg3tgkD2ZYQeIOUineCcM/b4nEkF+N/lc15DyyElHaqdZdh+blgej/QPkzHf5AUtB
Wx28VHXqmYiHDbFS/Ib67yWdGXN1K/K4Z8Jrctg9d2NIaDXZgIWCcbUdDoLyzIQ18f0LS05e0Y9+
CtiUPGa/N2CuWZargZ/RbbJOP7RZMkdQtw8OeWk9AV7a0FAFWUe2pjWR1TdkcQzOmRKUjEiUyPv2
3+5Z6TyFXXG7MdxYAeZ0ytNscbbZtRsBSuZDtN7IVodsPyNebG4LhljTEUN7u3Q7SEriOc3+Onar
ghzfz9pDgM2Eh53Sn5/+0HVVq2s5wd0l4pSwKtjSWLW5g4BcwbtWwd87fN1iz5fJdpaRA/4C7Ugi
9cPN1C3nCcjQ+IDm7WVhdnrAyoB1BTInzJg+81ydIVpgW3g13oAd9NVP4MEzGe5KpJzXhshv41VC
an8yZ66RsHiKv/OC1qr5917HXb3GLftIAJCuYRuCqlP9J1ye4OvkRF+viNFtvdLNhmoh5eH/1TCP
SueHss7HongRH+gcvTFDNzsBp28nWA7JMP4THdV9kcdJZf/1MJyvLVkflfWqlh8C0v3ntr6jSMxC
1464OWDIzML5K2nU6tE8ZpRv47OImZ/R4YI28vyKouzN4p4PoxBBGA2FA2UlVnzncSVrWe9BMti+
oqyCU5yl3zkuLjJ93Oa2ijYnfmQEuHhf4/F4Lx0Vzu+m8xd64pG/IsV8U6thwRnVP+0nznQ+8bht
Dd/4rxMa6ot9H1mzmQyqt7yMqSiwlVlVOFAMt1BxPGxg6ylk4b6MSmH/LY/4+A1Rsj8U40v9by1J
Xjo94N5AF8PkwJAqLi3WMfyhWwAjVVTIZnAkqQ4eplj62C7ObhNtffZIqBuy3HPhYxxLHkpJmhn3
CyTc8eOG+W1qgbnr1kdbUydD4lUKAy2KDZ0J8oksvOy5qQhu6saaSTGrIu99lQBISF4FRezhRgId
T9qpYBD6J5QRX8gWYioIcGk+9s2nZXntxQNwTi9Z90hDXb1+Vc75EdPb3n5C2TOxVFabQjQWEAi6
WtaWEVEpn043iDqHlmQqIDCLUbi0ascS6ZCy8bnQM6ORz2XRLzMVErFvx8NCLdL7PcGbhEcFtl7r
FMGoJI4RI3yZNSCOTwCDeBrJ4fhW73XV7ZIQ5b3/o/LIxWxe2M0qvokPYcBO6mER8T1hImBwqSJN
IZ86IlwQTrhEGCHwe4Ns/2eV2u5VtidLRlIt6+2MZhOY68+024kI4RnCzaZ6zuxQMch4ZJFTJv9l
L59NZ1vmJJcpl1vAPSMw3+iTxXFx1S5VRC5vr8jJs24Kn9zpYBnQBbWBQtKo+qIt7FwZCN1NZg7U
bwMgi31zKQ/IZm2zKFSi2jOuUp6oPRRNCTtByDW9xzSwG3g2nUkEnoMRVRqeF5d2w+9ZAc/i++sd
yqH4xK1XAbQVpQPSGnY7i9eZlCfIt02sWoFsbQPS2EypI+8b7dJ99pgTvaNIYZ30yQleghFU2/OU
BtrN51rAuJEgYkxhFNYydpAoLHkqCXyDgPD7W0mrhc+LUpxKCO/twrPZ3tcLo/2/6O9M2VahIls6
CSyaKCAE7Wt/pthdPO/6hrK0j9Dt3KQtAIb1WZTmOVn+dvx787lSiW7w7qY7yRVGmHd8OjoblLim
8v8NEvi+gopLrtkPTx4k9wiQwJoYs0+Op/cLe1m2UsKpkyeUoKu7ojIaDmkz3cjpB2ZrJBDahZhi
GblUvY6wsXX+63etJZWk52cE42FS1U8liuUaiOLNcr05osfj5IZzT4w92eEWrlZ79KzVASg0R8FH
AtPRAroK8JgAw41NIIx36XO9xGTp2IP+5Nb+u9iXlNNTQok0F008uA4yAbxIrED5F+iSApE/jBxs
PfOmFC4m4fffdrKGRRwNBkZxc/xtmxkxCvP69a7UUbJ9SveEFzFs4PkAWQkvBroYPeLAzm7N4zw9
KcG/7vE1bZmVhqqdDgUalLZd6bL79omOMKQBL/34PVtXi2hWLLUaKQ48cnHZ31rytrlIv3Z2YwzN
vdwwYdNLYAggiHbjEgp2ctAZs1+hko+usI9eJ3XZEqjxVGPDZQYaJYfjWiVkCpEiEzKrToEYRy0t
Epn2IoOJ/pbYWbRxEdaXinFo7t9Gd1R6avoQEYf4Nt/NWmTXMmsbnOBg5Fl6hJQnacfojkVIRdMm
PyM4fkeSNtL3rFd0den+LilPDgCnkM3tenbO2RFUqm8xjQ3rBoaRyAT7ePtyO71SGbC/YiA2G8sL
1fIg6t1Kkcym/6xeuJPexaBzwg9K0fYweRtbGKanOiIMXVJO2LSL6wA9UyrEEV/cnW/LW8UTX81c
b4Tb6e1e2LOc3saovykW9/C9U9wPAoQfdDBnvTxzhU6ew3CicIH2Gk0uUHJXWNpHnDdId7xz8C7i
5+TtD5X9FFo6zgbWP5Y04M+bxqKimL6aMo3BQkuWmQEaGZMzT/hW1o+FSPPiPXZNAWyc5S9HkWPs
OncbVwa4hfXBBNB+6QehbhojoNCAOTKbeQfeytNUFdEMDah9WRCgK/AJn5EFMXQxLqh/IXuK+CPT
5XEmb858f+MV/ZuMoh99MYpJMom05nLrulXL1CS4WBjXJRO2IPIg+L9+9FuIUwveN2djTXctpsiS
p/HjrVvH5pnREEI1CjgO+beccMKyT2ZScAQm8SjJOJ9Mb7HPjmExBJMlcurp6ecXUWjItr5JquXy
euZPHU1i6pdeEmvGgR4bGuAi5i/5sSS8UG2ZIdx5gJKQU68KvtVuK2QXlXn04Z2l1Tj/iJe1/fel
qPKgd3vgvKY6J62WEryk94s+sehymn71IgBIhhcNN35pbXzFHlEv+HEwfRdY0/Wf293lA3u2jC8r
jA7faJraPXJu5TPRIj2sUgzIKU6XMSSvPeTSU0BdFkQQt+8/V+lMRwKlRDFRMUHBbyNoauCuZ3zf
1ltHMODAq14QDBfTYmE3/GSFImrZ4tKqGbLClsgu/R26sH5ILlI3Z5XIdXHIvgtiSrdDKiwRczqa
+GyHrdt5iPdUnGVyX+FespZ4ooeyxkTYOjazY2pvjXp8mVGQhaLwrwk8Xm7UEeySSS/AKIKZwNgB
ZpkkYEBHlp2YLVbDwU8jCRFEEO6SqtZkVdK3n8eWJbE0JXOAn2Wzu34Z7oO21WMH//RCfmQKM61r
yTuvcCIIP/DDRprPxKEoyMHPu5zVEBMzbLk4h7hdz/jqqlcLq+ZD++iY0x8J9xr48CkvvuiIbg7q
p755XXkaDyQtRAtggEIzDJu2v9EZkCYzyOSFz+8daoaVI8JN7gkC9EhornqvZB7RJfjL9l2IUByR
ngwYkj2f3wpyP4uNxECXWewuM1Rlx5bpYQd37XPpHAdiakHbwh9JAxZhEQWoAR3FxT4Bra7HoOv1
md6NK7wfoyKZN886amAcDUqiffREM9WXDF0g4awpOP7hvTQhhlb70t4gDq8qfHq8J04GvbVKgZLh
iazJ8zeZ5jmuQUXv2uv/s9htOnXDi/n2ULssgn/B4uFsRLbwfQr6dg1qOkwkQLcDnoFUng3rVr7D
k5iyFJc0ZUGAbPjJM4ByjsDa2qWA4bvcU8/ujiKgmtfopWi1GQZEDtv6Ex+i5UZ2bx+D5UFJlrzs
GBSHgtk0RDM4fOc2WtqN3ABE4v+STcP8SdJ4x8epoUFC/VIijViCOtly0pwY7leR2v5xJIXU+hez
3bqvQLn2SMQFzMugwUwif61kG/5S7eARAiLF/l4/ewMqfdaEVvyNEibfRcnkcfdyjoe+Utu5fUDy
kXM8G8nZkMYkYRvpDe1ayO+/rOjHuSqrpkWSE18O8McOsnfk5J/OXDIGihGyCqiFBzAn92/lQrp1
0zEk3hDG838IRjBgPNhgC00wmUNsF+vhGmsciKopPyrdPVcGf1XKbGymeZSUJuhYG4vIcIwsCHBf
9ERuLmlFRLcTQJGIYsmSnWbavKEnzaH+ztXAfua0uEoawOEnvfLSy1IxAXYF388mySp6U6hyQdvL
4EveWUGvQu8M+YGpEnbbji/L2ovO9WuOTz6BI6HQ8jpHzLi1FuEAH1D/6mBOZ9Uwfk6ZJ835M18m
hFEcCiS1OXgrxFyzoSMmP+tOdwfhcfn8EWfmbOHtpCrE7Sp9dsB36LEcNGIFb6rt9/oswkGQ10qS
JxK2GF0ETjFPEv5VrSmDVka7IYyCTfh1SqQc1XjdMgr3zzTvowbbxNUlFerQ7pO4P2weYFgdQtdp
96CYB4FYtNimSyNaeLtMeZnzud6Tt2Mpondv26cgGsUrbR8eSNuy8b/fS7hbAhBD8lQkIarp1msN
TC3JDxTTnpCQ9UYq7rtsSMNWUElNKHVzqm12vhZW+g90g1xWxAtFjyu/Kbn14s97uMJEmISwUx4l
JhgGxLdWygmiuR3iaU4hsAquzjRhkNGPBAcdDWgLcciyE7rtu4nwp+Hy255xyISDrmHbLEknx0cA
3aSsRuKexmFotjbTMhFbDFJFPsT4sjqPDYXFzc+zAVem8Qg8DuLeFGyFelidGRVdXRlcy3fdPf0x
cFrSGP56UccWugxjmn62w8RpvlwQO7+F50dbKy61Et1AgTj+S8VFfQJu9vKzhsqRYf5UIIkaejb8
SRNZmXmv/KK5jW3aWy0u5+q3Fu8vpIH8VN3XuoFCYEl/mnW+DoMIjRbBUoWDnO4Vn3ZZ6/+sLIDT
DKq3vq/M4pZmw/kq+SgoNOJODFly/HU59sWbc0tzYio7W5Qig9O2R2QViiEo0rWtX5AQEsnuPZxY
GVgvKbtxbWiCR4C5YsdqrHBL438Ut1zxHtR4II5PW+vklKAD0OE+hWqmePAlYYHcIt7NDb9hQkKM
XL7T8btKX5GTLVfAC2I8bpCHqj7/sc0slJDAxjws6ayUVz0wZ8h6Tm/1/K+dj3MNb3G0mWNPJq9g
WE4DAKOs5SG5cI2LbbsPShgtMU8BBmC+vRYfQxz2l715cMKIaoUq/dM+4Xh1WC+aoHfZZrL4yPFq
GHkD/O/Sc0XkGLNA8LXD26ncfXOUT6YeJ8bai05/u6Zss4OCr4vMU+6fWUD8cOqhdGNutHwJJ9MF
EYUnPODYcBVZMASVBfyg+TK6U0ECpAs0ybvp0TUhfHtbAgChzbhtmg0/cPNjlitG9hdmLkYhUKtM
fugIfi9jp9WRoG5/szCFbcVoXEVF7FB1gX2SeaPdc+1BeAJL+4poAVnx7m0eQDJkC810lCxFs3Pr
kzBf288oo5Zn68BNqpCEF1jPA6zGt84tBEUnVdoT316b0nNie9X+FDMj6V/qh3Uebd2qfmzAGpvE
snvpPtc45vZxC+WxOtx0R+IuNpJK5isgrwEn/4jTovswqfzIcZWGjxID4pk4LLH2Wtnh/u8vzPp3
zpj/4Nfu4yg89on/U74Oqq2yOoJ6wrfUF5TiL5yjFEF9Eh7lY4eyDMLft9xF+2Fqyu5QhUWqJ4Ma
RkiTvGhwPeFbmMO4LW2DKVBobgAY7NYT3X5Ld/KJyrjSKqzG97V0uQG3JwFxyjB+iynfAeF9gge/
LJcqLutmOBYHATvE5wJSfUJPhcoxIeTAMjAXcdH/95JA/VAq2hvNtKbzQD0kuunTEU005vn9Kar9
nFGQKHyJwQbDG/exN/13hdyp6NomicQZGjVeiPwcbx/WGFm2ssHFnOSyRdws7gJeVbg594nAD5fa
neUZVbFNlXya+egvWk76mwxJnxWeChFZXbYnT9uRicq81QyZsxQX6z0mAIHGCTGJx8I+XRwcJh7X
TKwpwRmHbmpjSDuiJ/8f9iDOdjcZ8VjjS9xDqgz1yVt6RfTrdhjJh62YsrStQW7oMvkCwNd4f41V
aXif+thepuO4yzO0+6Ixl9UUjAanFCVi2+kGlA2dgljHzoEKfSYamYBrDF368+c0TIgpRuwYopO7
+R5T2ZOjZMVcgrpN2l2Nn0z9MPvs63yaIZ+qTSgJAzHnd+U7lPBU+KQZXm4qv4ZFf+YDMK8TaleC
fHavvAZIkVKPObY+Bnw3OxmaQC+PLnjx2xHTxFpyMamLhTPjtLmMoO+8TBgxKT02Dseei5yC1CKL
kYlZ5TbH9eJd2WU+rawPmkSQRf5HT9/q5337q6O5lZR9IBQ9HszD5KhddBPOORKn0hnw7BrUKR+2
DmkONUbXUF1bH2uvS3Qa2Bgm+Y17WEbbJHVZUE0adVeNaCKghqejtqANtfTc7HDJmigR6IGvBnyQ
WzoVbArJ5tyJuoKk7LGi/w3X9ac0I7OVLxsojFP3fmCZRzQC3fz22pB4dERMDQuc+ftnalpPoCTs
5ocorCypVVpTXE3wF82u9R+CRY8Bdm2pe2mau9IpTivn8BUD7gjAiQFz78kKobQo/kZ/B1yojzgd
sITb9pDe4HVRKaR0KTHSpsTN8gPuCGNftLrsB38LupaxJTTxhNPLkJyTOa+lyt8KvgGlQ9nZ4M2w
GzozTFYdoU7sqtyHaqXnS1vW4Xf0iWqFjz1fZ0q+/TurabesScYYR6O7cy1mQ08YJqckiRuxpcPi
kbSyyoJJoxxXb1sFIyGGJ6LRNRhPAjNygnDblQrMWDXjGzld4jwDY82ZyW8i/giK061rFktyUoLC
fgi//PCZZNbbEZw2wOiNQ19u3yVTY881zRZGc2daNL940s6V1WfTDFGDc79MVJHMaCZcYURrkTzL
0xfZI7e7ivWZi4Bfw5CgyUKT5z/VgtrHuNH+0gHxl2KltSafv63Yf5jjriiVtJZd21q2hzzXOHrJ
Cq2hvMEpwbZuH4hvghujI+lICKz6NETkatmjLXvZ3q2ceuxIhBYX5VFusbi4vdhxLkK4Q77rQy/Y
3YJuBAdOAfoDSu3lwbXH1JImI2Ly7+cK235SzkYEuX351vLp7VqZ6k0Ra0Vx6CBvAC1uiGzgVo8v
aHZA09dB2STH8D4gW7lafkEe6uCafmmcrWUUcYa4cVEgLAk30NQO3H4VitBGfIKoAVwwzPgxGP99
UQPATHoDn/e24nOUDUejIxOHewEdjMebowlcqMVgPz2Q+7V5KxRQZphMENH7VNVGV+O+Ks5Asmmu
L82qwVKnuDVNEuCufhOMj6rylillPcRFWH5XUXJL805aleFG47Z9KafW1VXzsrHZgxZmF7xGFj04
CiHaYXABDc/kc5wDIS4R/yWVbjzCkQJaY0iSk8gXvjDDV26pvQHFSyXnca0Nqfc+GxzR+8DHAvec
g2fyemRF9D6+sxtHkj6Ej4x8Kq7iS3BqA+0nC+daHwrz1Xx3di69bu/ySH2IKRZ16EkH05fPD5Tp
u3HAF5P3WCoKLqoI4DGMk81/Y/TQyltVK3/xx83Qrcnu6vUXuLPHNYD10Ap4TuKy4GksdPZnGMCX
VOq//O5DkDz+MOxb3rQKpiLZg5lNy4EpxyYqpeBzlQF1VRXNmFWK2Un+Gl/qllgNFSL4mHMOIY/2
JGU2Ng1s0B5zxbpUK1jQQVG42dpRtx8XoOoqQZI6aTIHDNxvT9R+CEKVou5gulVAk+YUmrm5Qkm3
WKv/OJSLpD7poq5yuFV3n4Dqv+jnq5pTj+N6adJ4Hrawi9YUBbgxDmtuqV4QH7NSLUZIIiwjQGv7
AV11pTy6J8wb45je05o1er5lJxWxvUS6AyWXKH7bVh2OsDSGDHlX1oFRTQRNy715MXM6JmIoPG9M
Xe8/DAnWr9AoSv73BwwEdtKG1lsrPv7oE4w9/8vU44XOpNRxswPe4cXxydVWgq2LplwV0uhk46Pe
KUd97s3VntqAMhDYcW0aRvimvIBch/nGMFScz4RkgBH9LBLr+aRliYgbgEyXfkYhDzTlZBKZ2JlD
xozs7emxnOi6oqso5/VweBe5LRZnM97fxqv0RGgxtKTu+q0eEragtha/x2osVbkAtmnkv2XfJiK0
Jg9gaImfZdgSa8q1PPAjDx3esopRVpf2Sxa/3lsvYxRuE13KbGtrqFlATOFLQbGUEDoGXXgMdmKg
M7pERN6v0aeOXtyjEqaslrrqshmjVCx3qA6ywNSYk/uArLvZ/609bGHfTZ5nBnbg9cdBa/rFUQHN
3gV26C0Dbl6elb48sHlQ92sqrWJ9hOur+KjtjPHy6/r4M04ZFKGE7CvmAcnCrfmRKzuvRRUNU7Cw
qx9LjOJ9VrxYaMRtNYtOlVtEochdTbOtX9EWQ4f/MyQxJWqsn9pCofEewrE7Hy2LB9eryd2DodcX
jNPBbmsYetXCbpf8ewBCsujr54j6Vk93xOFBZawRZP38EL5L0E8QXtvNc+8eoyzRfzw4F94LPsrs
N7MpUB3/RAY2YNSvNDoswuR8W8UAzSKyiLSBA9pGd5eYtdzpcc4M/WZl5fPy8uSrat7/EgLTBxZ1
dw3XU142LdwfyMKWMmseAUxpYGCjrV19/4ZmOkVzT17Dp/1rtD8pU+eI6chQbprh8WIP+glg762j
+g5ho6IHkLfGnv09HS+kqaTgBWrUhOSF4AHkwxXe83xp0deZSQuDGSM+EhEmzZ2BBPmfh1JRv8nV
pwTl4RsUyAPcMW6f6cPGyzel3WZMHScp3qexDuIWZdrGPCrOsRq0F+b5Y6cA+XBghU6nT6p+WtJI
CeLso3obH3Hldrtn4hjdBP7ASVjwF/1KqU7YO8GXfOWuleUjQgo7rMRtfCmlwGd8ETRPWlgoIiQ6
sR7Xv93+GqtBtJnW9qD70wY6MKSkmnhxWFIOFRZyzQWSX/qTZBnSGiK0l6VscE0bFCl9wr40iwDT
lU7whAWbTreML99EGz2tRgCX+BYrvVcGMn8ZTCJIAYXXaMicFuUeFXcQOuSyk7X54bavo4zsgM7r
VYwtmJgqZfHOzrHBl0fbMvV3sI/Hg2XWa6GBQJn0T8ERKig50/e3RMpPLlTkakngTlzyijL7ANQU
KKWuMbKqekP542ftXJCl0xoA2hRe5PKXzrD701FaxT6msiQ20cp5GQkcgJlJCtMy9TBybqzrt4mw
fnAPOZus6wfZKkeeNTDbSDhDZypcg+GtUV4z8gqT4IYeHGbLd8j8nonrKeYednoy67FHj3MohgF3
JaRP7u7ZoYjJKCNKUMMwpB6XtdkHIf9Y8SNQUV4CP80cwifIBAK9vLuCGS86QwPBjEmGxj9kYSq+
cX9M7LcOAAwfuq57PHjsX+nS4pSjv2Zec8DT5Q63X17cdN9sE44NCd+tWdhgfCy/tkF2tBRohoQt
aRZ4t0z41Z9t+bU4DxXN0lMKGVOeKZVt5RTANNZuv8gA4B2lyPrhx+pNgFoRTieeRScdubSlAuod
Zmt0awncpfAGahm7wiUnprqoXnQfv8uSduwYZz3Ytkr/jmfJp1EdHBckZ25j0XfSP7iTuDOrWZ4C
gTcDmqkEvP3oRyK1tnJZEsng+TGOhpRUdS2BMMzfQWiEsNYRHEf62FJ6HEhZ944b7OXQWCBi70im
7lqSitMa6qJQfpPPJR4ZcyvBZUb9/AkQgGGxOL32BJ+HaOnnRR3PUUsgqlBK1xH86TSFKHvTqtWY
gbwZo7A+gc+hP4vF6OZme63no/IX61waeHpeMf1jpm5jCUrT8zdD8X5THBVKZrF+qnsbYjG1SORT
jRQ6snv4WDE5DlVUYmVrO1PLYStsbYtVT/bdVAnhh3ok1qbiMRuJMJjljfdNLNNK2ObobUUfDrTz
vjGikMPkPmBu5GPxPkIVfl7g1cgAtalB30SQDreWCtANdNS9IukzIhNMNR1puwzIRtyTA9VlyVM6
dyX+8sAfoqQ2Z1hRUxDqVGX960DEGhwxtHYBJPAEAneZs0sDXL0eaEVaOlRSxitDZ84dJydcKXU9
10JMgIRRZz1U+BpKkr1tXK5o7anAkigUnWbL/O+tRic7vCrRrOk94jEFspGgyUIRoD80TKL7NnaT
VYKdgQS4XHOxlCJUxrm2qU1xELOCXFb3vbu4YYXue5znfdHs5YN/YfhoYwrPYzyyjArQeNT0hLzm
uhnTiseYAgIF7957ARRcJji7HwvkMEYxeXFG1SOG/RbMu5ZdOyCoT3J9BlbqWXFpx30rwCOR18Ap
72pu9pOuRZm4lw9+UbTyH1/9toHRY/ivXGUJ/E54CoutNiTFAh6O5us3oDiFLu4FMnkfliob2Syw
X6gNCawTH/AZ+/Lgo/JSTZL4aaZf2FB0zOAcFZEXP6M+BXswyQ16uUnMWT7iDYEfFLmLHPuIToVW
518BXD86Ulfzqkg7ALL6+mxPMyMjWNxk0kFgp9LJ72VQ9TnweuJDVZm/XuoaIjcK9OGmArqVm7dq
xuRiieYX+1zxh7rOIdQt/ni0kHNFH0UWzZPcGBBMAlndviyoVKkIPpC3OaUsmbhtKGdp8bdgDEW8
UbfABkdH1QvJNb61GruBjLMcQBaYz9dY+0paqA4uYPkYo2ElnIdlRVBeMVYpbCpho5MgUeOw4gYX
Eo0RViTBgoE/zMuvPuKbKdZQXyQNfQ26yph+szjkMUr9TUYkUNdZUxPOu1ck1pd9FOIWOMxcWFah
MR2K7hhqv+S7GxoGuWqL9qItxUU86a1zl6oMqfFthP4tH2i9tOamVbJ4s96r04WrDnIMV663qv3h
mBIj53HopGVf9X6EtqA+1gZJb5hXK6Rsh4mzEGHVBg8f5kpw/ypaa8h462gVwOHUDaWwMmj2I6Z5
MnzaQnNaOr1HBCwMYPULYlZ+oAjWidJ+FqLw5hpUQJwLykSYUHFpq09IDcgatMG/rIIkh3L42yhU
MuQ9+YF+UG+/AWGD8QRMEa9R/CiKqt7hOPjt3I2LT+vMo/lXqu5pe3t5lPktaabn2ahDn61wCerE
qKZJVa1srsQ952qAkUXsZmCobNV5sZF83Eyuh/Fr2fmtmf7jFMD8Ybg7HW5KNEWrDSphs3MK6XNL
A7hxOrZcHBtTLoH8dN2qJRKBM/4Orz8+LCH9pMs5ltl4IPLVlP4oGfSvABVfOaFiwxVX1H51OTeh
CmeZkreKaUnPGpTWEG2CSVHE2p77visaWn35kpI2H7D8srMECf87YJpVbuiv2S38BZBayjBKimZK
vRjNdjC4Scz7KLgKOrXHY+aq+qhtOnXtq4nsTsGCijTWtRcIq2bWLYxsczUzjn7nWpJxD1H2S1R7
8xT0vDLtFGBq9E017p3esENOwAqup6g7i1+qLze5ZwGlpzXcvrtnl3QXgab12FBVYwz/d0pPTXnl
MNGpjeFLQdSslT6pPmwd0LxcXmRWT70vYc85G8oAX+MWkRSe0o2xyp216fNh1r2G5D3rtzit4UsX
s+u36M0OxUaBvoHXOFVdVxmRheANpLPvC0j9AeW7W5LnhyV1qApmrWpK9yCcvCanxqWTBHo28PFm
FGJRUXZcy1yKgq7S3vJ2PiSI2U3zHPXTx7F9NdSHwpNossAyXo9ixns5s3GVWAANKqgL/NCUE17w
HxwS1t0UasDWNqwKwXcSK0phcxle2VyOTBlAIhC5HbC6mrLselMKtavQf/j0+/elztJ7BhezQ5iU
BQJeBM2gCdUrXgIeeOE6cnYMjBFS1mqp///ej14YipoE1WyP2IMbdOMNLkRXuowkGf1dvQ1h6H1q
TCt67z5iHblBFM7oaXkhP6ag97SOZyvmB+VrEhDXfGUNT9Tfqi/qnoS1kiBMqf46p0ABtvthvW2t
xB1SBXm/1mmTvUb3HCQje71nG7QjUuDjxeV/fFdOBHbclE+25cSMLEQqw+uH0+I3tz84IpUVIsu6
Eg/OOab80zZW7G6gf1PO6+T0F7hFc+9j9RDSdHgvgR/IfkBsY8u2RGhnKn04L1FKppi4Gfe2SCoo
BnmXlqrjINjh0uU2WjVBc+atVckWBfGy3WlVTumx19GJ+3v+JmkwcXUyeranSet23MunnmiCfzyP
+Ntt0cQbVL8WACnvEExm4zCnXhWK2SdmQLL/RHKi/HEqoW/kcfDCJtvTiJ4guCl1UdOaPZYp+taS
LYu7uiy3thAuEsARwcWsmxfUebMu6HJNtJGBeAdM/qrIOT6KG1g8tMZc+B5xbU71KBTJ9FnjYww1
8Upqd7csqsW4ZjC5KI3QkstMDgTDTi9tXook1/pu4Tk73vg7R6Bq+DL7oxIoFZJqxhwe5KZ2ZawE
/h4NH/3T1aJpMgH7D/jUiMu0VfWqq3eNwmp/V4eZWuuDQXLIC3XEBNE8PFA/zg7rvKXQ5MUsObTG
bEKMJ2kFn+0+dDT7RngQUIQA9CbUsF5ajfX6iS49jccN4pyfhK+GrOaQBotsEkchzLoPFVFnjiPB
Fkc7xKxPvuihoOjR9oJugjL0js0XkWSREJMs1eG6D1hZcYgb0nS0zRroMQJsnkYfC6d4LEc8Fdt6
F9VwsFV6S3EMyAlo9yat3tU/3K1q11v8dJV60ALjGiOSfzP/w1u4ZcZDvzs++uDlnd03PHYmh0Ls
oMY2WHhjiLT+nSmyTAHuwj8JL940AJh96maWlm6tV5TrQwEFOuwR4A2WtCBWlKLNX+aPnwFsws0V
bLiahwa2Kjqio1JvUIzKXQEzQOGhOWWCabDne7T7DUN2kUT1wGNg28MgSOIPvBjuCVOaJtk7KFJe
oprAv5JCWSjO2NSQUaUUOlbn3+1asol35ec4t7VFoD40anlU3rhbexLQtfyS+j+AvBX+prI9RqsY
EEXoxOpnF7+DXaX893aBFaqrnxkgfo1nmALuVgu7/H/7vBSwLvX54Zz+fIQsTt+EmsMPJSRRpiSA
kgsXFo6TUTbuPIqXho+ZPqWz5hDNKnT4JPlRLujeFHXSD2xi5QzdGj0mlo9HtdU5fEqj3kqOtS2H
hA54//wU1xTZKB+HpOzIN1x8CiJZFYl6Jy+LBIBiRBpgyS6ykUwYHum6283W+IrB3UocJP3GowJM
cMDXTYZ3m8GXUZzT2gbkVdotmZeQeMvGNyzZXHdO/D6a1w94uQMqvHCr2XpG41dHdGz+QnutoHud
qRzPkqsOoqwweyqjVcUnTnAf8w3u6588339gGfaDU5Bgmp22vt5v0I3XXMkOrhyptWsC+vwmP2GA
hlBANaRdqGGcwf7ozFCuEYfRDCfQ49yTJZ/xepHPXbyligxjLy/h1EaawjwxZXflbaOaWn1Hbsyb
jQ0a32eTfxGOUFPsOGaSZ7OFVdxQwljA5g+Zku0SFQ6oKF8ZvZdhvobvZQ9vK8bS8JlSaA2Xm1to
CX1SF9UcEW3/0sdD9B5oBuIjgD+naBl5B1gWX/N7WTvZ1qe1pIONRm+ErBAVoA+pj0GKs4YJewHI
kMoV5hMNZhIVWFmZXGIVEZ3ykwu9hfmOiB/O2sDYQjGaDcebEDWkn+dvwbWCpAePHJB6hjaHTB3p
d8ElmbLQqa0MlMFnYAIBynbiiS5yxTXbPNLGwHbr1GCljh+SwTlgf+zU0Xd0V63JSF5JXAdIO8Pp
1Vz/IjB20MrPaopFjaBICTsxARERZ52JX8jtGvCl/JnmM8XA38Nouy6rr3W0fzr5B6hOcd6p0pIa
VxsOAml7nVNd6rwdf19sTjS0va6WkaLoeBWt2K3Warz9RWXTilzONTi+PdIA0ieV59ey0WTkp0H8
h5kAXQST1cuEUzJlltCKaH/TwSWHnpkZjF7+YKy8cfDbs46vDiNvu4tSYpdpX6ffFeXSnhl197iO
/XE/55GHgKratmWCI4WcJRd/vqDrJUpjqmll/bOZ4sEDQ5/BKBjtd8dTYBq2+NPEHCmUretiK9dQ
Xs4kJ1Im6v/olUXyB/FeDSfKMjbJueQFkzRhCsZeRzMqaDpLMFEySMUdOtwthOAOARLTFRLWaI1/
5ttwZYemWWPVpstF2MW2kYhO2c60StfCWV44CUpaH10fJzgaq3dyB/0a4+96HhCkCiSQhYs/EBbR
r3YnQbGovkr4l0NvFEK+wFb2JnTZZC6Vc6mO97kHfud2dZdi5G/aovhHblcu5fgOwqvF3zYQuUq7
UeJ+jNaibL1VB/vJY9aukpZpIIgUvubzY2WfNmk+efSB18y+cX/+uELENnWt0qc40NqMfD3aAl+P
R4NX9rtKkVn3X23z4GEQ6DV/XuymAfX5xuZ+EVZHC+Hsj1MgzMyz4sccZOEkkMRv8GOkqTbAFpIu
0yyi7QtCtT3ksYDRCtEZ2t3i3WjQJXyHQqhcVJQT9foc344R9TrUV9Zrh5qs1g42HdwCte244qvi
A20JhHUXtG8ML0uRbc8hVtKQCi2U0+g273bZq26D1IrkUiK13NSQUUJEjg/+U1WkVP374YdlTA5n
tkkLQ7ojNY66ZPkJbZp9GC1YZYVsH6kjTdVdIcksl00QZvYP3+DRUuOCdnPCwXN+XlTZbnR/KRkG
UM8NfwiT0PqBPfQgP2Y2C+LpRJ+xM1mMfgj4cYb63o88rwDgUu7h2LAjpfxNSuLLBowBl1iM//Oi
aMbq5L4yTnX9wNoBtmuzwibPNKQcF8varRZNdwS0q0wqnUwf05ghhFw0/lcGXqEXnB1N35onI42R
LCjl/ec9dJEwh8Z0DhMH30KV91az6DPMkqsXAgnhrv0lbm8mXBdmjD5HyKptsGKLsG3hrd/tZx/2
j12MLpeDl4U9YOJVl5XBiLQ4p29RquXe2LhkCWY56dbGv5Z2Hi8sc3zQXC1kt5N6ECJnGXVkqQDs
nzQ76yLxlXE2uEMobuhFISWx03j6QGahFEFPABIPXaqLHuiUFtvR+DKE7lD1gubGeg1nVGPcIu0F
kJLIu+zZjqRETlD2i/tv0QF1VO1IdiJBxf3/bsF1EAmTABk9OQo9hYMM9/EWlsVwaaxGKK049bHP
X24icD7MzHqV/zexZ+HhyvnIIaVEapXVnIXa1PPVEhTkiby+poUOmToc5mfsoR95qeuWTKpBu+ef
EqVec9cXWprmeOSG39IEgzXChHFbfDDhmuS68MpdErfjxWuuk7zT7R4Jyz0q83PJE45TChyCCio+
Xi4Gg4s+rhnmqwAz+2Ukd8HYlhR2+jGPzMwCDf/xzybvuRoEGROpVa1lfvekAGD98OI6fOdQVz+e
9H97NifNho6IuWxtOtmwST4ZrDRvWQAf0/l5H5H59DscuoSrV1WI8VssqqlKD2USpZn+OhNqhWRV
V8LUtrRDCE4WSYwQOuZo/F7ujZOPfSqVcoIXnCN5xAT/G5XY+eumm/r/8nlm3Ti0U3iMCDsltU0V
efvj/C0zsmMsRPN+4NOrcPTEAp8DW8EduZGncNrUZ81M1P6/EFTzNGZcU5ITiTpoM7cMADcosBIT
m2Ak0bvABo10TDY3/Ca6NIdi1RiQHZydFqX7i2evjPpfQKh0xaKWb01wR1/aUj2cudmP5jM8Oy4h
eua+0ppeYhY8IGYdoJZM7VMFv5ufruY/OPqmnMcAxnYvy1yQDy8iV9dW5GfpYZTMN3R6wqUIGp8j
2kb0XIR6m1eZfWTTIg9HlqB/e3fKCsGAKa2mAEiy6qg1xC2GlwcY8g0miv3jkU1ylW0DGFnU8ATX
ZgHCSsT3z9MBK4AC3lKn14Yumn6IUrQffm0klLZI8sgihkvzYiHXETlHE2DpRIfw8j/IQ+Mp/4zy
4VsdiK9oX/VVhuKXJQmvsN6M5zus3RCoSirJhvUoTkH13itgsXKot3UxMDS4/cOdi8QQxfhPINRW
MERR4tLHBaLaTTyIE6pY6WpyTsPFwOiu4OaVb6BDem8dw3BnFXvLZPD0U7KvK8PPnsuUWt74+kBr
lt55yfQPGtfjn4ACeWKyKx3rjKZy2zpVZgDOm/DjX/FWH6d/31pS87yZgeujJmpbSqazttrFHMif
zFRREncICU2qhK73Yajs/W5HIEz4VcAyQKFkw/xtCsqmnU+9l2YQWrrmEvkvau0Fn2o29oSO9Orz
6tSwNBzWhQqZKj8jYM7Yob/pLNLsmwmF0u8rq/2pSswL6hStFcfDRuy7NPXnfdjSr79KU0aCrjz0
2wf6QH2+HEZGS3cHKNANBwH4m7pqSQKubo34qwg/l+rSJj9U5po4C2OMTYENh11/UlA03MRJ+aMN
1NRmNbx3ceMnZr8myv/6YjDECwcDNBfI5ZcaP3WSJK0e7nclZBl6IwgXFq8IMAVdtOXIFsB+mGFq
UOT+ELsoAh0quMZ03fZYl5tlNoFMgZ6SGDh3FL4jg/uzN2CROKqNvKlg29CpckBwYnYJ79sKUBB9
5MIXFks6GVadKU1lzfznAt42rtthGgnSAZ89APXUl12Q1cG2U1a51x6hsyvh5qcY81tXbrGlqhz1
5tJOcovHLLb8Tqn3V6p2CODLaDn7T+kgmAqAxds0J7a2vpcNtRzs5rhyvE3gr519G9opvrrrPUbm
kzxgsW7SyM8Kh8BMPVOJC7rX2bEOtXNd6idKLN/avCP0p0en9oLh6f/NtSAfjDFMLWn/r3yAgO/G
waxySpaZ7gr476ntAnojNT3TbRZ46gtlD+drH7rJkYMfQdPzXH5NHWY73PE1zNPr69GBzwBSfaA0
GVnPOGtP26w5e5eza6fJxSP4QzscT/oF9xji12nBqSrfgXgpHohhjb9LqYRT9FQM2ohfqh9jg9vK
6YiJ5GF6zaumLY/hVxBFptOLKXpUasGIw8DxIGQ4d8ZpHnS37+rwhwXVZ/MH26BB6b43x7TCkmNL
HpHaZbKFH/elQFcKIg9tLjyBNieCEyXO7L1RU9Wv45eY2xcBtJbHZddMws/iRRmAol/yiwOzqfNx
0FwGLT0HmUZ6b1hcmiRPOipMR7foR6V6rXtHYM/32qcs2seFy3B4yYl5X1iFU2CBi+5fhIqGncjt
VeckVhQsvrZmTxFLVN6YHyccaqB82+RLaBONjK9uF1WFB6+VyRxdcDZxFuViMB7KBWcuA+yI7Ktd
Nr/YWVyffhCbvJUfkq+q3cS2UD9NHeyfsf63mCTuuXzWapaDRv2HCoNAs1qYXr5TRPDqhyy9+75y
AlW+s/AyHtcubG0pKlCVdGpeBTQjErzXWOKDVNTEdguiWjuaByWeoG17tGxjZDpmT/uDoeCcsT/a
kqLwmhkla7pdVJrSaxykvrZautmEzwmb42GtKhMzMiBipu08F/Yx5cqNgZbx+7lcLc8u0vjLro6j
6E0rf9i1bHx4Jx1CCYkOW13rK5ca2Jgr9ttgk+Y5hl2rxj9c9nsCi8bqisecu+0n8G0ED+m611CO
aByJVgd5ob4SU92UmNKLpTFf3vcmoZ5XLV6/ifDskh2wb2tgYutvn3c6ksyl1rmXqMDVB3eMrYnj
sH0Jgqt5Or3sidfdZKDHYuRjX6sdR9VOj5uS7rvwBfn0OZH9GT4497GTFXIlSGjVZIGAOMjQVvSc
/BTg9pFI6/RdHkExUSH7LR3EPcj0/+ic0UrhshPI3pkOOIdXxnYeUNZkDw+hUKTopU8UO655t/S8
tGvUj0WCGVspmxGl/VZjQFSjWRaCHcOWWAun27XIvVSHv8COVvE6pE+0C3Z5Le3AZoSiUH0wlNg2
ZVSpP1WzMh7nDpRtLPO9DJDVY+eNPtHJ8g3DE14qBCQs5aeYOgzij9m5kApAONDbqMIzT5HGqpi+
MC60t5rlwyb1C8VDiFoSAdNfN7hOiflzz9gKE80REkBtNfpQ69zM9qp8sLh7kvViobjdWBPO790J
KUwZjGvXXfiYB7LaCOddPVzxNHD8qx0zevgGlmQigUsspipURH4aTHvs9NHYRD3Wo2q7vwxrIqsW
DKD0ouMerVgQK06Xex0ixIs8E0H7nhPePy/HS9hY4fWaoLZ+ABpy4AjtBgJXpzTz1zi1IqYkCxbY
l8KlHDpqm2DuFcg41/4r71Q22EdYq4pBvgpimyNpW05PiKBhsRRZ4N0GLFk9WvAnf7XqOEMTS7Ci
I5ArU/qhIhp0doFXOMXGtPHXYkIRCnoCHuLco4KobvFPRXw72WQRLvldfIA/SUHVZxNtjoW1Qr0M
G02f3lsCOBawtolUn+/wo6UyCgWWqgXkJaZB4jMgIkhCofDj3K/Xb+/zDeEeWIW3Sc1muJEVsACE
QDGHDExQktZwhZZJ2J5BkivSgi9O4u8wsfA3D68S/fet1414aF7sUQfR2oGj1BzPY/anMzieVzKJ
XE0xW40O/RHvBIFgaW0i/9iqCcdkulYO6JjEU8dkOH+XqclqLiTbxiSLP03fzmpHsT82DgtsVpqq
HNsozzRvzbwSl0CGpdg4jSpUVVbj+7EqmKQ1JoNiXl97GR0V+q2EcXQa1/gya/CdsCycGfSQP9w0
6s2fEzTFqwgNVkTNfXuyE8cyfBxUrw7QO+/ZKoZN0A1BEQlo4r4T3bL+UWW3KyDECI+9D/5uIs/B
lkEuP5pHupPL7d3MqfZkJJTZpUYJX8QyhOREZR1sJu7SzjQu8E+GID90/TZCKiGcFv+Q+Upi+5+V
aPmWCiX3o2oCVfkwgifaDH3Eot1e1bRDoz4vDGug2TLnVUXQSp2IvMW5BtO3erYFB2lboUGIeE8t
A0S+c8wwXXSZUKEi8FfUL9uw3w0CdMJmGJniBCmH/pwJlTavn42Zt1E7lz+lbj3EE6IcGgCfrKiC
kgZWkoIB7J9Jn8s+SE0MWBYzgg4zdxrt8Z3FzCVeje/b2QVODgo90A7D3hHo2xJB7diIvbuhVhhx
X8sZ83gN+we6U3LOkeN8vAosAIK9jXCNtLWZmwCn8EU8LN+3KoKpnxjBf1ElEoBajYYYazGaf6Ht
cwLnIH3LzKVMIi/g6FigMNMIXeco0kMMtg2evDKE0rEMDlwmDKPhg1nAJrSmXKxRsQ9TznlSaDdM
mBsWnIcULxb0wKsoYuc4rrdV7LLag/ufayttGPjyOgs0Df4H7Tb79gBpPD/MZo4mgJZzG212s3GA
nE3ulixun2QuEiJcJWTEwxesxv+a/zibdosNdy4H5JTsfNMGTyYuohQ+/k8bqrgDwP8sA9us4HJF
J8+Lut3NfgEfeJBTC4IHMS7Zy/z5roy9jshreLPVNMUkSsv9Y2mLwTnsJTjjdEVYXqW8WK4vD7lj
CtcXhzbWhKPnMhJTB4MTiZLdJJ6vgT2HH8xcTlKd5K68Xthkj0I0yMHZZx4ksQzdkdXj6YUXMP1z
qk/0ycFxm/NgOMLrU4LFZfjypFKmQJ8JeOswkH9/4asmT4LzXRnmAqjzjewk3Wt1bPWmP4KOzz9F
+SHtS8mIU1dXff4mVEZ/7I9NgP8BMZx7D58CT9SNoFN6kxgXBzPKlACVWGh8c/0c9bZ7CthjAf+c
5Ip+PuI09gwcpaab3dIalnDwcFB41rintSYv1HLP4gZ+FJ7T2wY5D9QZ7yILdgbG/7owMAfb7Jnf
KDIPxhUEcpagnPJIFXEjXhn2zLboxc6IKV1w4WEUR02KPdMPi6YUSShK8CJcXSFtsuQM6kPQjnlT
FbhLWlfGRmu8O01g+fNWnYpRjFHl4HZ3hBxz7NE/VDkV97NMe6jKrGV6ThZiOj8FGgam+OzAClK8
1wIWcw9s5GMTAsNTOI/Vn4X/ybgRleeoD0hh5DQ2MCd9E+sGIsm8tZeZvdC+eTBLpG9qerREGbik
cmiclK6pmIxwgTewMyJGstFNlXhzxaxERKfKI+XTTPyorivdNHPXNB30t7KRvY+6xNrJyFnUwXsq
gzYmZ19TDIRkEHpPoOUPEpu1byMe7tZIzWLtZVGXiQip8Jin6t6pb60EuSnMpiLsntFKtSDTXzt4
wvLr3nWv1b9quVFhi2mM8MZGH6914nbFP9zxLVReHoVTmlhrfnuAI8rfIAOuzGycdVOR6YXxUWGV
yS+bsTl3KIHA8xW6wqx4fW7GzMxvsTRKNHNbeT7ToKxAva+if9irqaXUwbyDF6Sd0hE68ZJ2rV+p
aD9B7rFHM3d7hF9zcwb1YcmBnT4fuvZepJeRvQMZkF70YJLbIUHqUnPCSjNADYD6ugUgjk+MebKi
/ACWeRtuEuJymdHkUKNcALfRkNYbgB4Xv0Tit+32AcDjczJ6mPXh943f/gCrXQ9lONyap7NukrHP
e6rj7euJiSi1VAtF5uoZ6ccnEWEA8n7td/gqA5Zpnhq+Oi7KfzFX7SQJg7RvjYIx8SFpEyQWDfbX
8rVF6nsFcbzLp9mHEYFRkaECwF2Wd6jNfaDSmbJziUYRKeE4xlqUT4rXe5G/N5G59a9yUVWp8CQ+
tHa9sZgn17k6aWXEqUOqlKkP41oBiSLHabKnAeb7hZARw6lzkFotDcFauq4ePbDOecRi4Q9Haw9n
cqbC3mDIjpGhtHbkIpx4K4ts7IyUl0y0yaM2ue5fRPISw2WJQBLF0wvS66r7NLgsfTfZb0TzeFih
EiDIHN1BFsuEZA3uka1zy9cw3A77dK7EwbH+EJMqdt9mEeR+Y3+OhRqgMuiMCyXJxObUHEoYpocK
KS0j+3yJ2z2iKTpyITjApQJucJJqdQZ93rmMusaiyeAp2Lkl/IzgLUDkEqARxX6CRJFwkjSfgExF
lbwPZAAnYxfkX+XSphaQYg5KoQFhVrMXsaVB/pyHEB1PVCkmnye4dqP6g9scVgZdvoh2sph8OwPI
cWBTJ+F7WPt5NK8ERjOsT3QDjjxMUYejT7OhGCxvFzo3La29ADkqfGCoVjE+3sKx3YXNLTKvwvkl
1321Z5PXaOokfBGYERy1o5heReh0uWErGbVuXMxjb5hYK/XkeyNdnF8b3A/gEQ32O4ygbdX5/h77
Z1BIXr2tprwOe7r/cN08mB2sMw8zmVY9IgRmJ214p+S9s42tPd42LX4MbM6pdlxRjTqSZkCMwzGt
ndqNhYf0LLf5qryOYMJdD1DpmJIC3eEiBfUfyGJDnQLUQc8nUhfDS3Mt9Y79mZrZ2iITsKUL4z3y
3z4ke7TthpCZzujDwIBu/ZbcZI7x1k9DYRHeiBqwzffj8Ju+M7QbUaH56gO99oqXzVsTN4y/6INC
yUk89bJ8vd5HpMx/mw3gwbI8ApeLNTPOBzM0RgZdRCbeLtY8Sa/F5m1DK4ay94noMaK1duwYfHIo
Zv683JrHjm2bMZY6YkRmuzSH/2/gQnDsyRlQlduPR+19BnjpfQX78k3a0Pm6n/CcON60hV5d25Um
qLP6WGJyjIHk2jpbsyFEvkIR+tBL+2mMXGwTuymopKL8L7pOJyL4tXAra1APFQ4Fn3mkOXjrW9Aa
/DkZrNhFD8r5tpg2TreBJBIQ/o5Am/81Yh760/AdrQqdgnfOa8VMrDa9BpJhrgevM99H1ineInmO
n3qM+lws/+zjTVBySk8TrqyEX0yTd4QM9vy3NV6xrIZ2nIjC8kej280CsacvoVcFhSPz/xRbfgZm
ZmDnxJuBAwMI0QF2/4RkIakXBxkZZNl/UT/ArOJ9jPaKLipkXmUL+Cu0Gi3nLI7oHZRrFIkdj31z
ykiB9OhwzNVZCzUnMOA8V4+D6gPcm/x/VsEkmmXIRsPPHJd0jBQEEYzdfxwC1cNe6+D8mEPTZmNv
Vqd9PeBG8Ml7bYs1U0yFOwACp8rJ7f51xU7sCYCERAGXBelqY7Fevr4Hfa/uudIFEJSbBntqOHaE
XRL0wRYq7dGxB9yep3annXdU/1B1GaNxg74Qtyz2TBgwmpCL9brQU1Tr0G8LO/MQAdYzq2N7zaM2
tmgpVyawvT0jHUqJu2yiTJ11nnAeKQrkIRiTfN5+/EQ8ntkI4UMzXRRrqQsMF8Tys/e/vViOkLxC
TXaqI+Fgsiop4N0CK2ycm34+RyrFXdqewxP+70OmMLbOHFrLkKzzKiBb9DcGj7+GeDznG1Ehyman
hm5Okwe/hZJ9Hlup0zOzFbODsBi7zB17kJOO54ioWet4E/GPDUHtaUhi+8BWJhvRPCrFWQYaaRQ6
t5Sl5UGK+kyUR2hy+0nwUmIygLjWn1uaksmR23c9DGtaD2I3g3iZ5uE55QVMvlxFvWwhLzPGs1Sv
7wEevUj11QVu8uZwO4LG3brQ+cuaEcIlIDD37G/TyeTYW1w2/rAO2HbHAMsvZ7tbisUXctZOwxqc
rmsEXvMmNzCGI+aGsJ3oftzWGdomWGgXpFVNQ1HRiEz5/jkeVsQ0/fm7ulUUrrE/qYKoUkWin+Kn
PyAXuAvk2ebpvJLu40A/V8eoRf6XvYAdokE26RLXh/r9GRytAC/xU4aMTsry1e4/soNuEmOgxjJn
H2VhSkujiJEZ+kXWUDd8d+4jH4xM4R/EPE/FlhixMbFQ70WnOi0oHWEr9lIDCJ1EXZRAAHzhADlr
3Dszcjs0doAimHEwhGOVwTb61IBc0UT7CDJHuEGeEUeA15FQL5ENkopdV6WA1aV9vKL53EVbjYvm
F7G7L9OW5zHFB7BskcWegTxlhcLRZnI28KUdOHYxDBEbdXY2z6jfuj6CaV2bn4F+lyXkFOzENRO1
N6CAE7Ms2+K1s34LtSp5LXcObErKy64lXQIqEtB9TxIJt6nGloVEtr+AZAMroEhdDq42qxl+6jj3
s5TBD64C5KFAchjAWur8hd5en3DyKcVCrKbWsvpXRIfzv/hI8PjHDg9C6cUsOGXqi17KsWFX5Oog
igCb13X4FuXkhtTlctdZeMj0gGZqowU1cgyOrmRnwfkxIKREJcEw2GIt1kx656kDXvsnphkbUQu1
djeXahoEKXoKeEz7QyDKQYn0ZPOd5mN3Vs/iVKoDtyNjX/qDoipQWt0cKqzmGVqfYcoHMaA/jUSm
XixT1MPPNY73Lkw+BQceFoqVA5ljHj7bj00mF+7imovfHW1A66kqA57wriqCfXEBtDVeoDk4MSfO
W1H4ZQXuh+DMIdPuTpaENT7WjeiePi/fk0spQ4iG31EVGIHMior4SLesfq1D0jtwp0TDfixLas2T
ENEexOBI75LxDQDfNnD8Srf/YnnvxzvGx/N9X5YqRrt6Inxpk/DgkvW0BAoynou7eYt4bliiCjTk
tG/32hd9rTvxTGg8DCIHQ6ZBUzaJcsK0nK8LiAD20nfGftGKn2kflYCQ5DMYcXQeuS67AZJYBcfZ
ImliF2MjNdb78XuU+CxvWvfHRfQUxTZlV+/VsaPLWPvMfTp3kSpf6nYupt3vuNwY0Yf8eSPwweEu
UHjhCotfY7AhgtFsG8KMYAMEcQqOhqkFaZNqBtpWxbAcQUlDz4Rd6nnxejVQTsMfYdV15mUl6gl1
p657cruixyBNFh18FcaJIDB3biyP1f54zQfOOJqpw04EzJDMB59CILHNfF7351altsB7UV4YP9HN
FTfWJDRfawTbU+EiOMxcTTv31+By/eCIGOUuTdcheeRrB/+HqI6sVwBhX0b9+7sdrfB6cBmqKyQa
WJhIDswxcYsJKeG0Kr0QdDsOjJdyGEFem1+5r8yV939ER3YyJ0JDDEI4C46a6rGl9PettVo6Btfu
NC0mzTnfBVtx/ZdqYjCsc+iK1VxKagt4aw1B+duZ+0E2BQJTmCw50sHl77xZ/bZJJBzpbB57XFyb
CjyMucAJAWCtWAIXn85LIcsrXm/wfoZfHNf4fuIC7OD5blZK6hAGT4ID+9C3uGjS/u+v2ZLpMegq
PdjSh4GU/WspbzMwEAFtqVl5L0SdvbSVZ0oGnsIGDIXPESvbkLOQ29R0+OZ4gm1bseJyoLV8ixR7
Y66HJrnmJW/w1Ne7AbL21nf+GpuW6zAsK5kuxCM7HIqNP58Z8m8qDC/q2fifRrB0NbkV1hlB1E4c
1CGHPRdsR7xRMARbtE4v3bmCRg5pA8lRY1aAPdcZTYOfpKGT5LC3MuTycAKCehsu2z8IUAWRQalP
4HYNpCeF/41If/RKV80bg0/PMCEu3MaPdFSpPEBgCzqoe8Oe0VJyfrQsnEDS4kQbeMf8ixm+kj67
ZztTO2HI2YVQ7oqoNoCxdJ3ZLTxRTNRXn5K7p9cwQmG1PuLi2jeLTXAZnIfNIi9TfqHvBArJWqfN
yuySLl6cX/yDSFI/G2XJxIaN1yeSv695O8Nzb548gT4XOiCcqZsTcaf4iIykS/QUPumVzR/CB9am
Rc5MxyyGgX7SL3yMeaGDx9Wlk2t5upp4M6S9OvZa96RLYDq5ThOZ0mYrjI+WT/2ZcUYdSSpMFMI3
XqgCFdRr7K4a+XfKmZ7InxmOHV3vjWK9mDL4NuPCeb+CNGGSVs61TZGj6obGS3ScjBJaPtBw0Do8
hZ4FyuyvtajxYvlvLO7HdnORQ8qtr/nmgLQIgClzFld5M/l0WyZulYE5g9jMsn/i6Hlyr0K2j8uq
pCEO5g9ExdpRkV4L/eUcChxspY6qpzDkrX3NUmz6geD990NcsNKi1f//gU+vBFkz/ZFg03DPITv+
LwjuoSOMHzRV8iBQtKDT4tjaXkkZhNi+cY/P/y3uYtihn5lyw6iI47ACKdlUh200SJ2uyNlnZH8e
Ig7N4wYq+0Loy0+zkl48W9qaIKIKktqF6axmkVTd9mb73xjGQddZvaolzPS6UeinDNzYCrbA3XDC
gR64RGSy1fsUMnvx6BoA1i0nQ9IottmySGBoc3CpJB+hPcfgDEF7yFCYozKRL0sU/Jts7iziYGqK
qIJFb/cMHaMz3+l+47tDZ/1syQk3NqhDDDRN0zyVm7zeLiiJe4lgYnaMVZ3IyNdr/E2fgla1SSWg
MVtIUAyc/sWMDecCxV2wULydso4UGdTOIP/Nhqh0s9XzKFxh1Ijoz2XX5AfF7XHp7m6Ne6/Z8X7S
8hgr9dQnNMXis7whxlt3luuzPRPKIjk7vlbz1b1M+ceNrFNu5H8Jbcok/wLSdi3lGypz/DAOBf8l
lKx8vG+8I8dhg4ATslxnIYzhazjKDdpP/owiPMU0l+9eAvNpAQ6terlXvu1NwhIPeElU4I4iN2Bo
nj98CD8VMdFCiY4uKjzd4GL2/mu+vcx0GUqPRSRZj0cIDQJ8F40ojr6+xtYh8U0rblfLUOOmYi9J
CnWABfVZMo42czrdByeqfkYdnkYZ+1uOZoqMg9nlBfYjK/yRFBZBbOHCDt3J0WQ+svjlREwtQdBZ
e+qTzvLkKjQWimzItVEtOYKsq5HE6GKqRjpSjgN6ClqLi3V/cB6eFsIy94gvXmAf8JQy/FWIXU58
s99VZcuxF6rLkLChO9aA83nlbKK3D6qD/CC5pA0XGGUwe2Ro3oT2F7eOUkkh1XlcjydMGLFBOk57
lsi+ODKnvxUq977DBxdpJDTW4MuAZiU8vbgamHK6rJn0v542hf+3eG8UvlXoPU65AqUBcDhSB9z4
gYrwy4a9XhajutN+K3y623yHxZb0awNEmzQ4P19Ua3b5it5hdkVomd3CPGDIAwgRpxvH53xMKGux
odsKWlMcbeEya0RNPKm++X61scEiJN+COsWmnMJYXyWNUjBeiYplWnqFzz2sLpg7//vcALCx7uXU
wnzFDz7pEffMj7jLmhw3ss41I0AQL3uSv3Wdj9McR4ZCbaJ+uHCDc8WCdAEmQIgDzLGJuIpe8NaZ
YzBUy/uSgRTijK5ZewM1ICfDo7bMDL5a/6xwcJn0JNGdQaT03DbaJ5kzG1KPb2PpO7qXrS2k7G3s
Wi9nSz1AVFZHdEdtvYKOoOxiOHgSoeeWioIVjAU93CiHsre7duLXpfFiC4bdL4OW/yAzZjJPI8BA
N/BH6YJuRGYwMXKZLNUt2MD7wjgCeXeK1MIDczBCiuZmC1xKHQU155IaYLtmNGUl1wg/s6F7wGeD
8xZJQYTw+z84fx/qCfQ1nTvkfOFuOuMT91DHq3B8cBd0KX6yYzpilldtU4Ntv1KRx5YM4BljnEdR
tEunA2tew5Q5DEZWkvSUvKmIF5IvOLd0eRbQTnUKOoJaCNwAh7vOodPs7IYjge3zkWFiOHOhw7tI
+yXfnCD+o037cArvvLbrRfPI89P4TaWjIBdXoG1PL2VeZbPBOUkB8cKC0bL03VLU4oSpMpiTooSE
3WxcKR699xPP+VWIFMVXCeQ3LdOBFeEZDOfKUgFq8xF+Y5Y5q7xP+1ybP9NqpZreevg7XaoA6qJ0
KQ/SZTqupLWC0BnAGc7zc42Q08pjBxcK7lmKieZgr9/29Q+tBy1XbQsDfcGkNc4kLENZJN80ql51
5w8HUSA8l2rKnRzz/JUYWl8THM1hBe9s+Xkmf3yu51SQJ0fQaDnykFSUqRW4FP48oto2/upiQsGn
AmHWhT+Z5FwOLtQHpjCCS0AwVnc+0O+mRCRKM8jYfVe3DRte5RndeXcECdGAWSkYeQJzLXiaPYhV
RXnYgYXgPSp53HurDQli3gEnM3lUa5Jgk0EKysbuWMAG13ZTEsUAEXZW6W7Jeuiw3C2W0CiJVwje
YdYf4U0idjVWxARi0JbCx2mVlWlNlFhBToqC/0ySBXyTZL0CkJWrCxMXjvxt+Uh0mKrIumZGaLaG
v1XJqa8pbwJXogAVxdlArFGbcYlLVUgk5JbUKWyaX3uywV4624IA2W7bnGY4iGaW0U9TwcHEj/ug
8vWUXfJUqaPLd6Y1beT2ZEy+z7a+TE/go1eLMdf20T39xQ4m2/M0X4G4fS54qN6pVWi5OtaFZ+oW
IDMOHYvpKbunSoiz/n98rNWL5Ei2YAUySK5deq1quROyaBKur5K9AilJlQbgNWL++wuh1qzP7ASl
WODV2wIswbQ/Eh6iS/63UDhgJN/dqbPTlSHvR+sxqfI55t0OEwnn4ORH3FqbIxmjWaqiJ9Qp166d
lgLZ6IBos6MW5vBnZoTAPK9BuWq0Yzo10sO6ZrdYeK3dC8DkfwR7wBSp2rzs9mhcprY6pOi1UsLf
GJ5klmkR0fRcvoCAQDHHuJ3fRb7KEtA8rVDI+YTFuN0coZv/UBBVWWtlnKJVxXrT4ni1dzNO+562
E8UktFU+FtdSLVOg3CEd1K/IGJxh2yxLZeoW23YdKCGb6vgZChWDx97W5Fvl+1goQ/U0BXGuhT0r
MSK22YvYyBPPE2zwX2jOyE1mHGlgfKFCfcLgz2b1Qu7TzqeDCHS+t52jHV2P1c6jsG7++ZfWMpDs
LQP+a7UZR3BA8HjCDAc7uWFm/ftxSbc8DT6w/JoNB9Q1VLI+zVoakXnsA5Khr+hg88d8nimePbDF
QxxJK1BDkkPxn2apLR0X9RAtpRWr/XqeEZqUflql+3arPgDkbEjvb4GeT6j5WZUVCFmtgWgj1sLD
cGFgJ2rzT8CRdLzrT5ZrBTwFSIjFyoXDiBUoX3VGMUsVTSAFntEn6PMYKW+sLv26XfoIjRo332gb
nWW8SS/u5QZrJxWwe52KexiBu5H9gpeayPk0Sam1sA4ZmsjTXmpE0no7mrfG275unSy20JCxp6/R
AOfCtehg6OONlfTDNeh6pp2E3DgHuBsQgZLauQtURB25cEcJ9e9JcGGlmtr1amD/Na5Ie+Nbc0qj
PZ/BEwODtyN6cnLzSwTp1JpjEE+BGmEjAPGUZxnXlHc/1n4svWkknXN4RvNdLkD9oEJ9P+Fqe21d
wSYbKSBnTPao9sc5qAdCCImafOezwcCGEj/WfIK7qIpGRd1n7/xwFWhlWqcOFuI9eC2/CyBS9B7a
5htoQL8UxEOma3NX5hVJ5rqrWu+e7C9uAzkQzMmpGc3YOk6JbTwIEjJvRNn05+QcyEimxgGFOZMn
EPspVD/fuFVwMrkMWPjS+cU3h45RXqma5h5txfYgl2Pzv5vbWeppWfq9TVsi16jCiUAdpIF5TLDq
GlMyvZxfK2XAlOL9rsgbrAhtz2j+HlPfl4jNqV3Oxi1+NLdadZunZjOju1mmzZRkeqr/ZjEoCVX1
Y+V1yTWbWuXdKkOI7sVkdS/Q3Lfk2w2N+jUTir0kZRqNG6dwdfYey+dafYSqJ17twnVWdJ+HsqjT
wL8EDTLiQQErFAIsofbJnUF2VJio2mlSwjG+V+dTpEvWVVXyRdTqNg2mOx/xtjRF1Rvjkw26If0R
6vKQ3bc8dXRbwvPT2EnkSNCz3vOC6hNOqHehP80fZFPECGjnyGAvFuG8CMOzoq06upKKoQPT/5CE
DMvlGmebajyPTwXJXQl7PjGFUUnM50t+gxD8j5mGtleqwfN0fpmrSOYQ74b48xJppKMKBVxyTaRn
vniej+PRHABb6z2YknwMexb+25AcV8o4+khGoobuzdvu58PbG51vT6mBefqlD6SN/RvVseviAeZA
NTrX5SLySjfQWBgSvuGKior+YY7dWgBRoSD+b/4wBw/tjzLjr5++um/3hDZ7EE46pqnj2wP7fGMu
o2qii1dIey/I3vl5uDuwWp+irNZSGLH2tlQbFmZbyz6SkmvIUHFN4JuNO4nAXcKuJRtT2Uigc8vX
nsu/xGj0XpJI7XgGNoFQ1/PouqMmu4doGUwZkKPerX19aZUQsv3/mKNmRaT4BrL20XTQiMdqRa78
d9/RQWr/ROfiH7cGOEhYVcPGA+LsspRBJXVOjY92jlHF/kI/4ADNELhK/FnZAX/HwTWySLn894Gl
EEuEvWnOhjWyzXB/9fHWdb9j+oD5jpmwUlCbdZJWj7imagwKoYw4RdI48m2hkGrA5HkDLz8hD3Tw
jnXhpJfJDMIe9aV1DrFegonjnNKi3m5bEifiMZ+ud9MV3zGNQSLtOqfk4XK1HaXesjI1k+5aph3u
5AudIwc6mYxY/XO0MjYOajIilteLAX3VXI1NmuytNuiKZyefM27BR9OJujx79ObKo/e0j2zJYQ/j
4DLFPEwap9+FOA0PcR9hXaXNHNmnkyoIOcaguXF8eJ5cIRDgCzSCIIKO5hIYp8TUNEtrJtwASUrX
XRXDa3YF1XrytaDFECnC58nTRRrMRdAyWy8B9JuAqeuhJMjPYF8HEUPm4Zp8iav+brK9RDwRj8hP
TdKFy/IsNgoAL1VdTpbZKFt4SluVnKR2fka3OsoGxv2HDNMBl/TgziDz0ltRQCkBIKh+gawIXVql
CkBZnCEUPjMO8vjxu9HmH83kkugdlrQDmU5tiKlS2Ch14+vMYlDVK22K1M/0gxQTTuBCtxD91J8K
tTmDKnsMFGH/SJrn3GjW3v6mdxpRg4qj4ubOueefIUH1rhvjaXyZXe4qoY6mbysmPIhnV462l/ZC
VFzBHGD0SYCyEldSGM4ogEdQxB5VgmL3tXB5O0zvQRxjItfX13zJWflKen0yHzs/SJJWMyxw9+YR
DAhv+rOf92b0y5TJKvRH1AzQMF414y5xyAPWkKxb4JuvrABNhfyKv7g9+cm9P29SyttbUiS0Cmbf
TkwYI6D2IU461xSHjBrvt0hP4rYNZBSaqq0CF0PLM0911oWIpoWwMfaN1H0twg9rCKq6OsrqSwO/
Wg0YNT1mu41w4mQ9FKG16heSo67ZMN3kPc48hDDI8YfAABkp1NewlHjcb9bnRgjkHBtm6P8IeXkp
7dv60RruuK8dkx95ATp+tk6FG3KizNGSknzW+BCYF2rzcpqcPKarP0Lm74NjCQs6p3z36OGprIv0
pEfJ7c7E64eaVDXLz+4ujxw4NJr3V8yPud+HCdWUWcpF9uZBQyCJaWHAqKW23FEE5P7lTfjVRb9i
+9z+6STtTzw1zKn8NFuCjPXHKqgNoF5fREw2ppvyv+TdFKunGb73TaI40WrVHixY5bbXE8mpJ5N+
KwOx9a8eQiEyFfkiQdV4EhtZgWAK7lRHBEsF/kZosmkuA/iBT/pOzjkX+d0E6ISdlowNyYodIByw
DpsO8jk3RTgk1UFaVhwIkIMAM/qsPut+OVW1wzTJlFOWTBMw8VoOb1hA75HeJfblUTC994LYEdNc
E5/1f6W64nT2nlelkfFyX6Qut3yqdn0vKqO9sPm7Sp5IKohTHDeL/xXA0Wb+kbMeIItggFCdnv6B
lexkb9mf9hchMbitZuoa1jxpmV54e3uSx6kAaUSi5ZIgKYsyQ9fzcLqyHpf/clH2qxJAfX6H7/3Y
sDsP4mJqiJQ90uiMZaOlhYDiPgeG0KvVe+AxqZZaTSveQ9kpuo8Wu7pzq2qxnq+eV96blnLUGgyA
ysaa0XNZZlZ8NIciZTu6fkm51AgcFdvpwqpVAoJGrN9o3f9zf++ASo5WUQUbKwqTyJZ0OTbJVqza
aRI38b9h4ExwPVXwbJInfcg/DiyF8XvrsfhBLdHcX9IxZY8kqeD0y2/ola7s0Xb9Rxb+ArSaDalp
HrnEVHQt3YRkn9oDOP1KBw6/5zhLBrp4meJHdMkRDMAwKugdHgtr0C2IoEdsrTUez+Utk2ChQ/N4
EMNxK8/JcCB7zQZAH9MAHnRNnuAcwe91sAFHM0U/RcNxoT6rLMcC8UkXyewmubYa8vqcNYdtvR4Y
KcavAnF70ddbjvrF0B6Ofb/3g/gRLA+Rj42si3QP6XgBqrh1xi8Jql24IqlpjJHy8yrU6fQ3bmmN
2nmdjINuPt0ClVVAahJERCoR67fblOmkpsxoWtfudh01O2Oc+W7xQINT9vkwPSOppoMPnOPa5t9A
3z8yhF6/N6BK/XdX6LzmRIG6U7IR71yUffwGoT/ay3zFBKnKWh0KjzKeWRia6OKem80NVAGFOK5Y
d5JVbnbqtJ8VUU7EMs87gYed+avUhQAVFh5yQZsDlrT6iyrPp4oZ4tUh9rCSYoZdp9Q2krH/bZO4
vQa0lVV7C8caou5YbM5TVLxccS4gYtCNMHARCCBx9rIVfW/0UKPeBzF6m5w+Iv932ejXGSJwF6YE
ZbwNHZ5/e/1VMKItMHTpE6z0GP/sj4O3sbvJpWcUbBAXw9QwDNrhvzBtvs02qTJhdVD5iQLCRMXz
9rkekiJ50aEdSBXcYIvWy8mNbhLVcB+tfPKIwnX14bpMYAaU+5r9l+WiH0dAOPHomA1g2xMDaAXk
AbliSM3bkUUiLikczVLfDRlP8PmglHdpxNzoY3Qxgi/QhbTa39v/wu9W4D3AJvqefOL+qGRlbb4K
1vsu0vGr0VfFMxNtOp30VSjH0/W8EqrknJ1MyunP3ZFjsPvxieRmfcAxDH0xdwMBwUR4bOFXwHSt
cRmi+ofCckzxgC5eDfbW7zyNoamxBZMNdLEeg1mVOFg7EabalXdyCtnTYVHIYXgcKSC3EdavXG2t
Ge/2c45ad8zLKJqENnFAsyAdiyEJPmzAXTbePVJuPrSwJbLO5dDCK3Z+De567q57oYf+wp7ThqPn
0Phx6IM+cTFh/SyAfwJW7sEBEcpX9hSUZPN2Zi2fI7b2yg7flpP+M7pCzKVKZXbjEosrrz34ogTz
dC+9hY+JzhSPoej45YdCieVo/JPUpMuHU6zrmtxmt7AQ52A3Zr9UPTQix+Zhr/GzidQazNy0cAfZ
IgfNeGGeZTBxXXatQvoBRDoIGop1/UeEaeTuzdE4ew+WNVFtRW7spmqozStp2NUSfDwW6DsarM5C
zh10E2HQCOIgLBCbGSpxQjVMeFW3ZDXs9g5UPINw2qFEhErXnPZmeo5P5ZQHvq1KIhsu+i3SCdku
QakGzitdzVCSqSri/aZIz4Nf5fNxreXxnVy0oBAhxqJW19u92Ruazkwq2QYBp1m/mGGZhutvS5QK
GdGhWx8sC+3I9eXAW7bIu1auOXE2hR1tr6enAvq8BUw04n+YeVzj9lyFSKrnbE1IFDP3oT47gsVB
dCCnfWJs4o+752FdcAS6nLjrWbPo+d47KvE35tbzYn2JefRdmqKiSpu9jXcG4BTHb0HW+uQlxCPM
HrSv9rSra5MXEybmxtBvM6sHtyLvZsl5ZHSary/8kOC3/B9GkqoaRMPQ80PNhw0O/GJEH5gvLpZC
clTchARxOkv+BHzPc//51cZkYf5dF+fxcTY2Pl9s9Zq9w/aCD3kD5t9D/es3G1MR2cMjgRvEl7p6
RrBnoI+7i6YO86IN7eM8RpbWe59xrLqCcsUKYCXecU12vbXyCeKQn7Nf78Zy59E/A5V0Hp3/D4hy
Z0zHm6C3pR24VgseQ2yu5tOWdnQE6fWubJGVaMeqvVA/4rpAD6pCYxgOudCyd2CG4bAo6exniBC9
+JUTOoTOmXW+1+13vtKfJh/wy8oCD2gz1QG5um6huc95HzCsZR24U1GhL4FP+Jc5Pd4xTSX32Q/g
G67Q9Y31vpyCQOGmXhCLl1JYI0ocnLiJv7+ZDsgZNQuXS7081mIVQHBUtQKxsNF3UWQL1tVZgaeb
GfHq4atL8SPXkutBYVcEsu5iyq6MTIdVdhogZjBwXb0KGaSMwbStdL7esOxjxpuyMwjCKmWqb00j
RJ6b5Q+/47QrHAQyMpA927JRV9uBzgthFvTGfTs3Z/jx31OjL48lcmS+5Dw78M9LKTi0DtITFd1Q
qxF2UKCAhdAQ9jomw4aTuiD/nx/jNKaZZvJ5+q70RjoJCiXyhPi6x7vXsJdcnWDpCe7oFhQ5seEL
YSpAkisl8D8ZcjbQrusrw2TurOUyjgeUiwGIz/mQuBXVi3xwnwMyeND1ZpG1m7UwndlOEF2r9b99
JaXccnrBYr1oiirYXuS0WfoP/AzcUNdxXRMCmyRzxN9ikb+Gm6zggcF9LkZAii+6/2cDV/SHJ+OB
jBB+VHGV/hNTkWknIUwWjmJLSczJJGo/sWa5UBc9gteeT4PUpw7yRt/0O+Fiz3MQD60+fcwzPK2Z
eyV6oPgMEH8WrMtUNz46Z/64mo672MTFKtMyJx4Fnl5U4qiaRA9BzQiKggO3eLeYzg8OsEUYh8WC
/USDJTszRvdfi/26ooEx89FFdEBMyQSs2Wh3yA1ogiO5VWWhYtEqg3/HRIn3h4UvGORJswIa1HXG
RDOUYohrwIyYpjXrF9mcHFw4Reiux6CfHaus0ggr5fJbOh7Mw2eBGC16Wsj5XUnoC0Qmu06pxuu8
oaLM2RYBCKsv9Me/zIcbZTAJIpY+Xy23s4uUotLHsZKxjeBusPoNRa24Mg5J7SfbeYSk76+C4CT4
vinKnswG82iSFRiFT5TjTpgraj/6amX3IiAG100tXilYZkP2iCmi4zojxD/Lnl4Kov2ZxS/hvMBC
8lO55r/GU3cBRAkxmHZM76QAqOqaPnvDC8NShfADMpNjCgPYa96rz7fZqXRs+LYbq4cleev8mxaL
w8OQP7/ncJfzKSgTu0QVqS6HxqTj1xQRenUYb1inznsYtNIjbIBjJNJoju+2B81N592bqM6G8pBp
Md1NTHJ0QzPD1HzRissWwSHMiOj4VdIhrKQM23lrlraE0JdxDdCpCK1UL9TZ0jxK1TJjqeZmm3y3
hEWHPXcpPfgfReYpBHp6sAGnpIYHgJqs30JR1PdOApa/Kh+AGIm6bVzULdbFOEEImkg7zARANyHB
gPoMuO6At+ffioJLk2eZwTkkfTAUqZUi/pfRmWfuj1u+f7FgLcT1ybYD4/qLRJ07QmV3wlyjwPDW
lcALFL8INe//U6MFoN4AkhVmhwMhkkrTbcz70PUQieEtTFt9iT+k/PhdHGwcVZcnXHHH8Mp7ZWoW
L5VNCVv9hDZ+JCKgLOYNG51ljZOqV3uXADQ5exvvY59fcDgFIJMSxu9BAF7hPq0Xsux69nEWaefg
VdXTg/8YtSZ9K5etGnDHkENhg15CO6454kEQU/5SGqEvknENQts7iU2rOJ2pPQUdK4YsguqvSloX
tMNYCJWj+CtQfSMrpvLIhBRTJwu50u3qoiHSkhEpX34lgKLHVSK5RqO1w3QEcXhfZYJoW9AiVQbG
xJEA4wsCuySKcuwc8vdi8EdBeKVADHMaU+85dSEZNySAR69cVa5VECZZ/PmsepDe2u5MMJcM1j2s
pcVnPzY7lJbKW807z4x75HASzpgKc3R8mT8YKirwyVpWBL/6/VUa7UzipFQQIyzIBlKEnUPNws1x
JZme4GFvqFqqu5J1QS43FnxCAsAWTA3V6oCGlGylLXWeIrCq9T+TRzO8sICxHMBXXJUt+7cc59UX
95IY7cLENfnRceil8Mr9XoeA9YdPn1MJdzYECPpsSc8WncgdnU/DMJRGI1BBLBAzdFnALqTRC4j8
lgsDYLGSsie68tl9uLUwSfK9hQlBh5jlq0TwcIHNjt3wfO8Ida3nZl8y91Ja3MYMBdogJN+c90R6
vY0daUSrw3xekCc6VPQR139FcweA7rZrtYMhccS2DW0mzuhFJZW24V2FC7AkBZPsdSnaeal20kOn
UAco4H+7/QgeyTbzEw44T1TPj4eXmRqtUXCQERZ5PmCJhWCSbbNT3wRpIuvqG41J3v2AJKPqVo2L
D3smfgkURbknElBLqUNGg28b3FLP54DwKvcRXE+XvHjUiSA9syFXMS33XcgCfN8hAFbo25vJPtKQ
3az4yATpO7dZb3RUg4yqt7ultUcgQwozPU0An6H1fpFFxGVZY8DMGc5A823TA1s0Um1Hux38YaUg
MesTLsGRKA0z7uW6FmRs/MU8OBeMkcPIlcOD49Cg+nG9WjjdO3Nvj4HW2KZ8Cw1hniTZAruemSE3
bOGXCwwuDjVlbeykquAQjBEEQ4AgBydu6n69Evd0VCJaRu75R0V3Ur5aX8GMRkrbt/xT2KpYdxkF
MhUxRUp3OCzmYdJXe/lYa++J/H6MJUZ1xAtsny3zRmbOxpLRIvzdO4IoBMAvuuI3vQ1xy9JlQQ0w
5IeudDBnaazcuTAJl+zBpZb+YwDJI4CsoXKqATWU4DoBqKegIqmA+80eQXEwPNGWYN4Ol0a36JBl
TlOkEE7HgBeTPMDezqO8wmiDAICppETMar76RYeI0pNSrr3dYFGhvj4S8t36jsNKmPEpKWvIq6Bo
XyDjxPVTY7EeZnJCBGfXeNPG+V1FNBauwWU7EbW4+Q4mwI8OEFWlbSgDU9k7joh90hPV3vbXNqP9
rSmmhdNmgO9X2qlcakU8NCblDh+6+OM9x+4+rsRXrLeNTI6jYE04N/wFLc5HZHni8aVreUtlzHvf
Kdbvkokk1B13r3/67nR31VfpmmUb2shzAXMhgGc0XBT0l8zsPswxXl0wX/rDTPnfYD4AdbFNH5fl
xw3fTHzpKm4TEt720W9jL4/c37m/uojTvmiDrkpHTC4w5V0c95Mf6zPOX63DUjel9Zer3SJWUUHs
nLvCxv8ljYA4lAJwa+hv5ReQJvmPhyeEHwF5e+1jFGamzthnVkjzji4SuRo59BsauS3pWTPbUni0
UImgQUq4nCkAI8V4EiOxrLRAD44bpx7MQKahqTKgZwR8Q1tnqJQizkucbReHAaDPl7vdlMHjWr6s
KftsrliTzWw3+hfPLx7LvsPO7iYIBXNMGbHC2YJFhPThv/70gquuiie8KQDWdpueHsNicWOS3IMs
YySmTOzJq9VuapRbxZnfX0nlEkh+UYmw1cTRK5vxF4ZezRHrc+Z8QASgdwzQ6iEdhEP4Jw/d2QIB
cAsoN2S5y57M3U3yZ/td/3nXGDZFtOUkif+G5TmQLUEAxT9q5rGkTssLdhqXcEVSppBDuLzMa9JE
xzdIhT023B0VQ0PWS/ZN6yKjJx3i68SKrzJsrTbk460Y7ojn6JNTI8lRge/mBrWbQEnIOHMCNTHJ
X7n+QKc6ohGzZcPJ4PtZdQ2VesIoO+4mcYZDKNlqQF+kWS38JqN7LacjR6pxV0rgkCj+CBZn6FQF
RoLToi/jT2IgIs0mDC9xZYxtw4WoE7rAG8EvDFrN0udz243uo55b6s+jTapJx1OLJLaB/5+oGNah
YD9ryDck78pph1OVdm9p+TTshazPYqCwOK0W0C54YX3jjNfSAPIKeVQg4fJhSxDeN1z+hOrPrbEA
HMnJ8gpERpfT1MioqUIchC1skh0pPqW7FdWDiqXQbTa87otmCXdY4YWYVHUT0+eNN6Jp8+TvzIMo
PQnhHFMG54nxc1gLvzuRZgJmttWTnByCK7vcFMJ523uHYS5M84ti2m6vKAodhTS/qqSqSm0tZ4OX
2d+0x/y3Nxkm5SPxwl1W6oAiFptG0qLi38Slx9KoptYXiee0RX0gqw2+DWWpk88eKZJDREscTIMr
IIMskpE1VaXmew1iLDPt+wqHaqKmjDymlAxCDuRlr2aoSGFV6J9faunBFJ5oYouwqgcStfGkirhY
qpUd8oLb/aQ1IdKT7PkIOVsz6rU+2oFMLQfttvh9Jpqb2D8aVx+MzU7iSXdz1d8fBH9YG6Ue2sSb
Mx2XPJy3/VyXWji5bYUXoPCDQuoACyBeh8PUoAakJ+4RDig2Xfs1TQIfJSfQpoXFBqlUrS4nl0Ml
WW/SSnuWtev4cXaef0A8b1jTbJilRjO/qaY7YAQRIuM0qMdL+W693HH0H+Iwopa9xJLeHhA6+tJy
LtxcN1BlO8MrE4jjbhNbPT2JiE3rvVdWaY40Q9Tg+Dr9ccV67pZhw6pSDKbShWxOCMVKxU0YOlzI
1FpFUYETEdsLvy7iR/P8QOTnO/ukYxl+f5MZnY4MCEFFxPpqrOWDMPqiehzp/V6SJALrLcG8KYYA
0id9p7uLcvSWzuO8iFh3TBfEgfPqFTzr/GedQ3uuGObLSNgASDAdHhJ2TDRjrhdjap7S8+xTfrGu
zca7z607J9xlF//QRde7ZZZAUDTfNMw/0FoLazK0eNoI+xsh+Lt+kJmdAOON/zwO6h7aIM2m6Ddv
xEN4b+78+TaAuG9+P24hlVYqOafGeMD7bMlovWskOoMNeOTHT517Nhpynv0WN1qt9E/qCZYvYUZd
GFNVDpBj2SD1hvQhKnbeZ9NQ8oFG2hesLpsPqt7CzZS8TRMQTdGOQpqeuaxw+EEQZwk2mUP9RxvH
MD9B4VQEkQ1bpPTR7s7xKqzNhCG42pz3sb+QrJfu77iN3wS/gsAFatleQBHLcejUseJ8nzjDv6dI
+yZEOGYdD1OT6+sy0kzXLfjokgHY3zM4sHU6mj9Ze7YeCmMmjwaPhg1ZnrAnqGd1fspnjudCfrkk
OM4+mX3R7Z+KBXR/glX6aIsEj+lO+OUX4Gbmw+Ff6mZrwaNn9l3NgRaRpCweg19qEenmwQyoU7xt
4sEvyISK4370q9JrPZm6UzHuIauwKrwhRVuQBU68s4wv0kJzg/2oEA8nc1+Yz3XSRNjiQR9lLlb+
+JZzwe3sZ1pA2NOGrg6LSSgKFlPNFTW2YmXcRrPZ+odasbKTdOMmdbrFlxbpfm70X3y9riNKHek0
OU8JwB32q7RtC6kOlbjVowTcQxqn8j/O3L3fwdky1Pr2UJ7liy2j89PIKmH4xqk0wt7x5pDlQkVc
gbB4UQG/J53Hbf03Dqo+c6wFhCijB/pcnbYdALM9xOvx1ajng34c8HSz3+ofROG+aibKeNMZ3zdM
Ty7By05lVsTeUclf+7XlDqhJGUsMMW7Hk7ugvnKHIu/FZhm2fAADKcSYt5V8YNGUt0qxWb95bMxT
l/F7oPZUtxdRwdQ3pDBMuygvnrKbcXvgeJ7av5EE/XejFoNW79FI7eTblh56WdcZweruVi/vC52R
s9xmR+PSaZjSWN1wMaR5dfhy4sZF743Icpkj3BLlPUgsjEjFsfGIiSP8M7WQRxQF4HRj7/h+nyb6
qPhndbnTMBLtlspz5jWyEoxP01P61xTq+O6gXUvAfkioEeAUecv5G4a3EApWoobDGzS8MIf74mjs
B19hZi/+MMFQdZEJdlc7LYzfVxPR6hb/Tq2yHivaSzexlefSmsg5OZt79Fvk0DUQyF0cMdbYslgY
tBnCUcSy/buRpl2rqsxDfBDb97lcmv504fc6cPax2Qw/jghXmdKXaKIaTx1Q9n7JXo9efU37Gsx+
rY7BoD6YQaY3P82CuVnVSK9NBf6f+HBR8Bcx+rIcBcpV7bzAgwCygrKQziBdoanRRlJAYuVbgewS
lagGvkFIU6YW+9Z5SZttbRFt/wmW1arMMxUAVym2u9gYnLBzBqK3px2/7I0TF/p0+hViubM6FnhZ
apSUZl4yW0YGByHiWIYtOKL4EzXoNv+g19rxDvxUu3gExpAdr0sX6DGWZJ5xrrdysBvbT7jGUpny
RjNN4R/ML0doY+iuijrd7r8bnuog2kN5gnjv1d6bHKyQXrBbNrtz23hxG1ESpXAbKBmYb7zsU6aE
hDrfBVFnB4lBf25Vep005QtHwevLVdTiq85ZSmDmPpi6AleRYmWAstwaPqMTKjEcJZAOWA0KCA64
ODoJ7CH1J9RQR7vk0GkonY1nLpW4XqbKJcuVIoUAP9Bf97L7ckA4jdUSulKAakWu7qr9wnKMOkn/
m6g9Q2xmTcEGyckpWbubBaSIxwEWsB2qNdHA6g76IfkQXMgh/tQsPnsLl5MIEHThq9WB/LnM300C
YVJvd5Sj0VFlE+NfDa+QE4//blThSQu2eDVkzRGCD1EZg45IcidTgIGd9rgyHOtKd/vjUjUo9Ipb
lUv3xjjdK5LBZXArpOqSs1cM7A1HIaL9rF9KxVHO9XUyGkDCEq7j4XC0h0D9yi8n0hDIDB4wqm6x
HGiMm1Dqsrj/4QJ5OG1wxT/CXEsHGj424u6+g7QKsuCSwEicr1eMsywEutNt3dEMODHDN+SO+F5H
WOyYBVYKhImhXPfr4kIKM2/+M1VtJigXd81iUyWk4vf4nPWW8GeMSKA+ozcKXptiIRdxv00ny526
cuzCdzdDojLvE6iUHgYttCD68jtkUM0koiJ7sLiHx9TLIzVKe4Nmlmrgo7S6oc+Kec8t2Dx2pYxU
nRdFZMymdTLDEENyfDh2Sc2Qj9KzKUPiL2i3cW/dkTgW6cXGmxVb0dMC8NITau4TWMlcG6i25LEp
p/6kUu29to/nXAsEtZvrRBC+fZ5SVA6vIvIec60nMpR4x31PO4KoZO4UeyPb76FM+Rbjn4gPwRmX
2OeS7vorIhNVYLtPp/BWlF6KR+zMfPbWeTyESjoVIbMRrLvdPCKiuFHkOuVKcF49t93MVH6+IRnk
1+ie5zlJtu6zOPg6kyr6S5MdgYgybp3xhYPx61jXDOrTxzxa6b/7aqMz3+j4SdAXUGdpLrUwcF0L
qlD0Gq/CdKR2H/+WMSrmtYgsVUxqz0IFNo3aZvRQAtpUXZnsOg86DeW4IjPK1KH/QB8WzYG4zq6f
6j+gBmnV/8Y/EtyovbrjEGKbv37wW6fpGCkUXKn3PGDcHorVs/+d++MqHPnKr92karbiXueqkjp7
W8/R/QPmAa6Wr07xbGYT/+tdsfzEDgCS54wYJuO/OHop9KE5itmOE8L/M3yvFKYF2kX/T8K3CJxV
a9sjRwh7z0o4w+de/wTSazYuR6wCsd3l60fcFGSX7GWZ3MAPbJppwmLsTLcgm4XTWdorGq3ZMbyN
FwwLbHFlApeGrUyL9sf7yOoPcoTxu4SUN/l/QiIamTTzl90ESfKnHXX1mQKrYsbv2JbSELXYKvQU
N0iNAXtgxeCb+9r5GX/Hzga9X8D4VUIpSqE4d0fyc618xHv1KvjJmu0ZBedbnqZsiJTQ9IThyID2
Duf4O7qFhCq/zSvCNlOW6d+2I8pjtGnosr3vSvDwEtL7Fbqtu6veIW6r2aAC+KIIrOpWeYHJ1iNB
6IjqfacbaYJbz7lW5D4dyCyc70LRg6QGPt6eURtu5nneIZLDcB9wmZ5aWApF6AnTJKptZ8W7DH5P
IVsElgVI42iJ9oQvy7mLrbaU0KHwxE5g/rIUapn/Fm+PVXiBkYvj9EqTuZGrGtyHJNSYfeHel7qd
o90Nbkacay31Xjmpw4z5qavWFgeOK4WElwCnuCSMHd2gWxSJIhfh6Zb5YLuJjG+4bDkZI5WwUA+x
/zhRZp72fK+KnZeKfOEWD769z/wtkuMDewRgD6jjXdTATbZsUUB9GeG5NoJZiWB8ny6p+wCg2px7
oRDnNlVJ0/bbC/I2f3ODVqr8LQ8QfjtQfQcJka2aKIpqIAIXhaxzztmVxfZWKixEhOZCB0GOK9FE
z1drcO64b+m2ROpkoXiWBbWHHZAoUdpbNq56m0/Jcb/WjQy1qoQ+9RpiP8AYnHNmq2rxjGj2eOW+
32A/afaJk1eITt8U5B7dG57/kAt/62cXkz98kdHC0s2g1vjSjDxpaizcgupLECmNVaI0+ZAEUzwL
hsvOLziHLh65A5DlWwl0O42Zio3JQEw+ib3GTE49yOvt8yeu2X0ZL7aVIcPfp5jn6+0cyOT6lV25
xE5nb+e3amZPNpWVoEie1kDuVI7Eiv4MzZ7CZei2SD/SDlGoU67WnSe5t8dHry2vDdnqJpYUJ+Bt
yNVJ6WBt3bhlxgOsNaXkj5NeMnNgWBwOnli1nVej0sDsdjHOXQvl0od9ONJqrWthMfw6mJy/2emy
Q+MpK3PjyNrIxP8Rx5kX3eaHgxAXz8yJ72pLsu/Rq1VK53VVLwtzrXurMawyvmRJML8Yi6Zquy6/
KrTqqZc4R+PxYczba9R3GowQ0FenLQGm731mvKn6zLxbPQFIAgjTTcecFbkrXjUmu5oR6aO9JdkZ
De6s3jk/BdlCrbegxJebPi5nDTID5nOBUiGRRZdtirxw8rlmTvleBY5o+iOUe0WHpYwTPzmVtipT
QZmIvcdoqqht4dTzk8cbVK895u7rvVd2U8pn7mnFVkpO3DiNJXN7ovLbY+JzqitbmP1Y7AjZVg9s
QsID/UvGhfkjSrS5uBnTM5rZGeZReUV0LT2IDpGv/rdAVbg4vW75Qvr6e3FdHaEehSidU+Uo92mH
Te9eNIoJ5C5fS2JBzan0MCNOs0OPHfsA5F5EJVYoeXtg5KEd5f7ZS2+jKU/kBAKUrd49wihbrvxn
AEP+d4L4er26wKngfUZILrECUOGU+c4THQv7WVD6dryLCeyh/CfiVq/GWAH0jyWa4i+TBP8kkMiH
Moyob1zaHIpbR/bcAQTHQzPghUVUxtjM4rGxKSuoZnMKgMctqYfRkglAkGXcj6U5rh2Rdr+OqGMq
o+xOzZ0++798EIpywWQQHoW9iuNUK6VCoOl2mGA1Vkb9yM9SRozsXDZudl9LGHxJI2/GDqb4hq83
cFapIaA52k1YApnZw9wNuTob03bgxcrTfB2cU+8gP8VV99yVIoXtHhqoIHwwP+GCtccWT/NjcTfm
IA9ix0HbFvghp3G2DlL0jTdQ/lEsL+pBk9D3KWLP2LkCMc7xAZ5TmsWmHvEgpGWyJykSZy1V4M+q
oWNe+QjOpGxoknEeOehSHpkutMOjyj5FqU8kd7oA8yVAEv0oMZ+M9blp+wc4TtSTIltFnvq9rTzK
lAFuQKWklX77EI03O+D/brO3D/+Fd4CwWXdSEV+LE4S7WRj1NGeGozrCvbJ3qgpizYlNa1Um2ssx
fZdntEKmuHJcBTMxjGJSnfaxnPDKGseZhXWfOECir5EJ6DlsK/gDpvCafUDnBd3/UZ2FEIAUqAUh
kRtlwzcEUnJu2QhkKkWpUQfUY8UqOerpESfjfpn/WLAVmbGYmbq84xWmJZjqgIWsKlVSfzLxnz75
Swk8DH3Wl9iG6YR0EHeLBs5amkuHVenr93CampcYofDR+puQmeb1uc/Hugi4nWY4d4u9d7tqxb7c
0Pb6mKERSYaOREOnC2mcXm82DPRqJ4Swnu4YjT1vSMF4HZZEWlP38bWK4Vta0n8p0EvXG2Rm+mze
iWlgcZYlo8xirJD7RYfXLiaNuOxDMen3QrPVlVJxnE4ceVm3DEqIRO3YhymWT7c+fKtGItQtXQ7T
u8pn99Adcji1HV9Vw9ywzutcdej29CjZvCZ0jsWUAGaHN7Z4P/1IrIUiFOzvMVII6hYUY1aX1yj4
A2Yrx7CCqSpL7NT8GfXHSIb5gMAzhXUm5IxLNZv0M70tiSAGuGJTHMRlmCIRkE4oVSEHADeekv/z
61lRHOGtwO5LDqFa7YroXNPUt2rgjBlvE/UxSMNirgDnk0aAe3L8MsjCfU9FFQ2/VI0Un/lhxv6a
WoUsPcF9mSFbs4eLyNDZFF3wRGjQ6XFYYk87zLZyx34F4/2eamx1Mo/bbG0y1Mp/7a0Gq4QGY66e
LU7IKEf5wZK+HBQi2mSkEc2Y+J9Hz4NmiQ8JMAPtLcyqq0QmdaBhYR235LfuDVp5U9iMKb/YEArD
shDpCAUWCaxLtvXeNldQ8lNhEAZUnm888+lGCaEswY/P+Td+v4U20b9Omrq1RhwAGTtQAxIPqV91
TG/ELy0wYjRwVu63ki2LaY/FKsDaaY5984T47cRjZ/N3wjYcgixg0A+ejlZ9e8t8hQpL7od+fl/x
qnzAAoJ5VcV459kvnRGroyOHDFBy8KMxYYoagt/3edQF94s4v2PyFZLXi94Uway5RiZDlyDiwmCf
G0Sw3QPQF4zgkUZ0kxlLTv+yDHBtuZQg7pZyb0d3lTbDx9vj37A2QcHQlzYuIunIGIMNEF8FEerk
MPB3jr+RQuocHRo5E02ZMlYqKm0bAvq3fza9gYHMkTM//t+dk1sE0BY6cH7SqG5GpM3dfuJbbLw3
sVy3gyX46/cRq7j1F87ncZKZadCJRzxwRHgESO8aL2GXS8lF4mqXPutjXEhwbkQM+d6jrXzfR1se
X6BAhofQamp+NodzdMul62Dw+O5o/xIeVXGYvdderbtJ+nNR1W0jEdM4GOIHxvkPAzdH9iQlLc+L
bbfQst8fgGkSC3Dp1U6rBdDtDsKTVUVCZx/PxNvUYVjxqGAEFlqxyZTijz3TEXI/xIwoqNeNZbrL
/0L28NO9Ngd4CyH7a/Pj/LAmvqHKlinrWqObZQFTEZjj82Fg2/ET1sQSi667PR9HrA6OedtnJAKk
tqFUxNS8B6sO1LOXUsxHBlT4BDiB+RH1BvxrtnB9saz5aJKsjI5po0uJLFIPR7UaxT6jPo0hFhCX
0ee9/HAuKCa8J+4NnZ89vy0iCzUHx8Vxi/uMb7LnEqVNdFtGihdAzEEdbees9TOGWo7afh6YQvxr
Lj5xuwRRZmmYh43IxZKAII1pOAYgp4j5E8dlTWm8GrTPzcsb3ZkSpBrG02fK6WJxmJUKfubhuZJo
fxoE/P3VDm4WFCLxpZi/EN+13H4sgdoHtiW8wLoZ+E/nCViqYpZF+E+YwEvGjoVu5XBHZ/JfxjmQ
3No1jJgTF3xFfEOa+mPd3mzXQSZG5yRvGTmtYffCud1sG0TWbnk8YDIysrqiCp+95cl37JKVciuG
BPbtwe29V9V6oFF3DYN1HPQ5AqtkQ9scUPDWK/ogv+MGRpV5Y32Y322ZsaQ62x+JixHFgZgOhMCV
nlKYKBObkWMtuI+Wr7YinfFtav+QhMgTqjjT+O9Hiyn6QJ6L5AQq6iGkzPgrhUrF4qyVis8w7DLl
ZuW3l691Pm3sof6dcyxoPbzrmOMb1gBXoiCscC29K8sNBGR2xlC4FvQbANM5g4MNF2RdVBgkiR8W
/ooq8XOVJ5f79K1eB7oLEP0NNrgsP9eqRx7ZBOxwPoZ0w+kAQd1QF5Mjcn5p6SyZUMaD8SrKM7yX
5j7R8Fe1OS9K92rdk0aurFP3sN85yg084y+qH+rtPauC2LASiKhjNZHvqZ1OpFHVz2rme3+EAiku
gAmwd1sZv/rpYdp7snnBc+NyRMfZaZVBa1R/f2QbfjxaUMDVzSTvIfLRysE2Jh53Q1LN+lbjGveU
5Rl70mjbYHZb6txNJK4VowMMcztP0hknDuiVtPZeAVkd2rC6AocvjTZxohJfkDNY+iUeltQpRKtF
LXREzrILAuUEqQLu2RwT46srjottyDKYqSUiE9HjYDQWD4Anw4g3E/2r8pc7ER3W3j36adJPMgRn
vXu2NnB0R2Bj+ZesBSg2eR7lsDU0p+pa13kkmk4oJRe9xvIhNvx0Q25URG70EwSCYhx8aoLCoK8b
RZCIfDPDMwlGoodYXEdLsmSY2opkFyDXv6pCmdSqfmMczZzt2qn/agkN7o/tgEsH1bHySU+AYJSa
8IgAyrMPbYoEZj1IhfnlvR+oWZeXRcDQPf0hu56yQc1loQ+PhF8glnJwGv/VAa7BC8ALDGHZhXa0
Cn+0Y0TLRKS/vY3jrJPuONl1s8myhq/I+6oo/0qIXPRiBXoAd4MYcF89llhuTd5urLWh3MHulDjh
v8IWqbp61Q5aUhYK30dnmIQZZo021tc2ZQSgTDf5goXb6Njf6JAdFc7fSLZWR9CTbFIebSwNtbpn
X8kIcwN5vCNlckux3G9YTRkePbFA5bWk9z0/zdEkc7P5hWQFQqCOTIWnkMNh6U7EDk/auY0rHqCP
cm1SZLvcQfwh1dj+UMpJPf/E3Goyc/o6B9aWV2bbSgRVR5K+bSRMFM7g/QAbuhEMO/UYyhWwEfMw
79eppxGQabmE3tIoME1lofhJ9eMDdbLqVLoQbouxP+Vz7ERJyRZL52T/A68dZVzikXNG4y9HuzZi
p5p5rdYZEo6I+hm7H2PcoEqSeWUexSdHfTSak23S1SZPue0k4JaDTr/PUvoByDFY9fFHW/Y2f5lQ
xP6wiRFanYDrjYDCvn7fhHVVcwEFL7H8Ayf+fRqym3wDvokScDMM/ZtBmMOQKWOLURXkpEJeLhcC
nK39bhZ09KdMg9iLNtGQ0jlq/r85likJt6hqetDBNqDVhkvnasngP1RygRsUAHIaFtok6GIN2U9s
ArM/8Ty5uJF9hdaZmw9xaVQPEs97yQokqpj2HymdYsUhPedYNQtHHbe32RQ8YBVeBYAJAVNAUvaL
bzOa1/eb50o1T/AiEiqK1omOZuv2FuBY6vRgbFJ+fIR29v5euMI4wzm9DGGloq1rBqR2bPIL4yvS
G3t1835dc+pMhMwQnPGCpR8P4v6fF3KAMJp/1EP3UYvH31q2s9EC0tautvttKZD6XwD7FYRvJ0HG
9IlIfOHnBJybKub1MxMw5/ATSGrUgnzgj3xVv5e/h08xpf4V/0T3aq/cLwUWYR1ka6SF+bY2r2X1
bS3lgklUtcKh1yuwflHdg2KQekhRmOKEWsS+OFvXIbiQoGAr6g8G04GZ7Uaav9rmIx2HjXu6efEK
faXN5k5533jHpgANRqjdhzjxIYMzviTHHJuIEVRQvyxOde+PjMdXQluziM/P9sY2kqa3nWIALykC
BMaH09bwsmXBOIuXX05oHNleNxK/AoYvrRu9YzWux/FGX1hufjz99lla3dfn21HzQN+C5B3TS6ID
b/G824BA+c8d18gMIzQ3HLtX3WSHEdn1OuwNK3uN8eoj5PGeolPALVSrC2YCB1wwaG9g9U9Tjxje
JHelsrUsj+cO8u8cbWOIc5o0vZsks2N5sl6fnz/xNAPT3Watwlw38ps7v9RtfjFQ4gzAjOe6w/f+
L09zwyF1FgyssNrF8ya1c+blMkVxSLEwaU+BZkF6N8UNR+xlh2M8QPvs0iDg2cXv4H+cOgQF4Q9n
YqPQOyCpO+PGMsJpuDCCcu5Miq8Zo3IEcv3ycAEgw0w17cr2j7Wn6RBAyGJEtZeUqT9RJ4AGHPWw
/NUmBLNaEpsO9k4lHv5oo6niDf5DVxRHmlWG/IWRZVQdud4wEcTFBj9SQEwl7yEUKg+Qr9YP8Haz
VBbv9uf9EAvxqtQN2DaoMY2+PepRDdTEIROPJVJdmfsv5z/ToEjctYQA79Y8TZBhap+pQEKvKRXr
J8HrUIrTBdjiP5ZH4fk6RRIgZvgsKPmhUHkYHPzImvcir8InSKt4v2LrlsjPzK/ZSDvZOshVlGsG
XqEcZH+oBOY7B1qXUw9PeS1V/vGh9qu3omdyorigB0mSymJRar++B6Mu2W3ndRaj/4eOcJXhl14V
1JIcqIq5n5hjPK8sq5ahzkfHqsAJcOJ1sf2VA++EifZamGnkMruh3MXDt3gf9yVqAoJGgDOzS6Tj
CaGpOPA2Myi7eK8WnwWsW8ZzCE1lQ4fw6m/BMionyH0HQ533lsXy2qNQ0RDnlsTRfiFOvltQbrbT
lDJXpXq7EwHbV4eOQAb+zNeVe0lB3Q2LFvCpPzGfq6hEMGleS3mC51QvqjmZt8hruf4+Rk0D7DZT
qhFx8FkH1dmKd6a59tb1zlKYXcsH8Z8o346y9RZ+Xi2JbOhJAQU+soNEtWj2/1baG8oODfWVN+Dn
tDCDuvFWC+WamudIm2ut2PJ4Jagja/q2qOz0Z4J9mbj4+nYr9QRNPvFGHqwMKAWYIAEr0uTX6Wio
JWSV3UgSaRBQe8HFH16Az07/DZUKdelwJje67RL3t3h8Q0I/wDiGTib9iG57b+k5VeWs4J8xNt/V
5TAXKW29+D1JaS738yZlpq2TUvWwtDz2e0fkVqy9+HrcvlqUt496VrvIc+Gw1BQpafd4q5JdvZLd
iB0a4+EUN1dUSlICdLPpp21dRKSUUylSLjGh0F2MKFD2rCaFLiiOxJXail4+SOeP/Fjfz6NB6tTF
GHsTWZbPw5FT5nR2yE5B4QQnh9XV0LohjQUwyHEGrv4HhxvcZEtbX5UoPPlN1UhnYbNgJsq6VfqR
hSuWp9sQp21gklkNeTH5OrzYTbb3kyDcMoqIEGjq2j5qfq7+9Dp4bZyGOdYYOxlpwjPJZnB3NaPR
VqTEgQ3N4HPT2cUzlQJmBW1iCOO6PCNx71RbQuPvnfGTaeoU41jQXho6hIJNR7XClujwBBbmlfs2
NFqCSjq37O1n+kIVR2lzZefkZWfoJtuIF1/CX+SQJC4uHKNuTdbn9klBJIzbjWyElJPkLfAEJFwa
4SmriNshU0wYeSCSLlgxSoitue7aJddEY/lc+8cK++Mh7X7RHj11e/+uQ6XjHk2HG4BidWM53b0P
+3DGEKWeqShU5NoM5L40JF1IqVQ7nU6f2VG2yPLCiFUQCpI4l+X/Zs+7xmpirMiSdv9jr6Upo4ku
HEgZZWX/vPbnxX/PYCG3FDjyXz9D8klEJbXTy2ulLD5RVArL8EUl5VtgNxT9BvC1yCnNTia7X3za
cfVicEwuEwiw9UGT22o+wMBQEzs+SwnkKdFeETsCfhwP4HsqTlx80xeXS+aNJGbUX9epi873O8D+
XpcprSm1M815cgzYaNBeBV81qMLiOQP+/EFux7ah4TWet5PuMFV/c2lyt9MadhiHDVTYUeUMn+Jo
HiDcCg5yr7cPxJAu8L4inhgxlYcZsf5Wneenjj6C2sdHuD+jgYtP3+o2NyKtbmoKjZV089yrDO0u
kYDYfiRIUOaTeGU799gJFzclOlGkIdT2wHTjMWFFt+AnirFdY39fxdaG/1WlP/13vwmgHyV9QsOb
JQr2h2lshnLFjM8fXlxq35u2yKhB/DimWITQcV8GXIcPaMJ+quj2aQFcTz2AMhiFRlFKEhR6SR7O
RpAsIMKzu06a3BCfvlhiYwTjBae3DoWMAXOQMEXvc+nU9bLt0Ge85nKOBFJnIrnKcSiBAngAKAGe
qJ1kFIn8cFCxJDzcTYAdDso9XJpNhW0TZRkI9pMP9R3hYbbSXC1oiCpj/jCDvLyrB+VazFVBozcR
CSqaUDDJpRtNpjeD1xT7nNNjswu4U3j0SPxwTf2qmo6IhUEQPaTAiMHRtw23qjrWL5q3bZ+LzGZB
j1WCj4dZ/CIY6x3veIBt+HGJxRjq0ei6voVwG6Xm6Zs5R04Ygcgz2ismiFhM/H6MVTgdrJ8rardJ
9Yy3CxyFEkJGVMF56VEf93XdcHkfIORoID8u22npceY3Kbabej4fGOjBUUQs4R2ryEMQB4YHLQao
2l2LozMYJvPCCmpIe6E5iVcpXd3xCYe8D3shW6WfalZvheHxpsFJPL7e+frWGGD4ooA6yoDcgFeX
kw==
`protect end_protected
