`ifndef DEFINE_VH
`define DEFINE_VH
`define module_name gw_can_top
`define AHB
`define CAN_FD
`endif
